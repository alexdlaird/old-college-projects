<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-60.6657,9.25,25.5962,-50.214</PageViewport>
<gate>
<ID>2</ID>
<type>DE_TO</type>
<position>-11.5,8</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Not_Done</lparam></gate>
<gate>
<ID>3</ID>
<type>CC_PULSE</type>
<position>-42,-2.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>BA_ROM_4x4</type>
<position>-11.5,-2</position>
<input>
<ID>ADDRESS_0</ID>2 </input>
<input>
<ID>ADDRESS_1</ID>4 </input>
<input>
<ID>ADDRESS_2</ID>1 </input>
<input>
<ID>ADDRESS_3</ID>3 </input>
<output>
<ID>DATA_OUT_0</ID>17 </output>
<output>
<ID>DATA_OUT_1</ID>15 </output>
<output>
<ID>DATA_OUT_2</ID>14 </output>
<output>
<ID>DATA_OUT_3</ID>16 </output>
<input>
<ID>ENABLE_0</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam>
<lparam>Address:1 15</lparam>
<lparam>Address:2 10</lparam>
<lparam>Address:3 5</lparam>
<lparam>Address:4 7</lparam>
<lparam>Address:5 9</lparam>
<lparam>Address:6 2</lparam>
<lparam>Address:7 1</lparam>
<lparam>Address:8 4</lparam>
<lparam>Address:9 3</lparam>
<lparam>Address:10 2</lparam>
<lparam>Address:11 4</lparam>
<lparam>Address:12 7</lparam>
<lparam>Address:13 11</lparam>
<lparam>Address:14 14</lparam>
<lparam>Address:15 3</lparam></gate>
<gate>
<ID>5</ID>
<type>DA_FROM</type>
<position>-21.5,-31</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Not_Done</lparam></gate>
<gate>
<ID>6</ID>
<type>AE_REGISTER8</type>
<position>-22,-0.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<output>
<ID>OUT_1</ID>4 </output>
<output>
<ID>OUT_2</ID>1 </output>
<output>
<ID>OUT_3</ID>3 </output>
<output>
<ID>OUT_4</ID>10 </output>
<input>
<ID>clear</ID>9 </input>
<input>
<ID>clock</ID>12 </input>
<input>
<ID>count_enable</ID>11 </input>
<input>
<ID>count_up</ID>11 </input>
<input>
<ID>load</ID>8 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 16</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>-49,7</position>
<gparam>LABEL_TEXT 16 Number Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>-3.5,-1.5</position>
<gparam>LABEL_TEXT Double Click Rom</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>-6,-11.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>15 </input>
<input>
<ID>IN_2</ID>14 </input>
<input>
<ID>IN_3</ID>16 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>11</ID>
<type>FF_GND</type>
<position>-24.5,6.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>EE_VDD</type>
<position>-5.5,-0.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>14</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-15,-25.5</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>43 </input>
<input>
<ID>IN_2</ID>42 </input>
<input>
<ID>IN_3</ID>41 </input>
<input>
<ID>IN_B_0</ID>17 </input>
<input>
<ID>IN_B_1</ID>15 </input>
<input>
<ID>IN_B_2</ID>14 </input>
<input>
<ID>IN_B_3</ID>16 </input>
<output>
<ID>OUT_0</ID>33 </output>
<output>
<ID>OUT_1</ID>32 </output>
<output>
<ID>OUT_2</ID>31 </output>
<output>
<ID>OUT_3</ID>30 </output>
<input>
<ID>carry_in</ID>18 </input>
<output>
<ID>carry_out</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>-48.5,4</position>
<gparam>LABEL_TEXT  & Average</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>DE_TO</type>
<position>-37.5,-9.5</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Reset</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>-18.5,-48.5</position>
<gparam>LABEL_TEXT Average is just 1st 4 bits</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>DA_FROM</type>
<position>-23.5,-9</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Reset</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>-35,-20</position>
<gparam>LABEL_TEXT 8bit Full Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>AE_SMALL_INVERTER</type>
<position>-16.5,6</position>
<input>
<ID>IN_0</ID>10 </input>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>22</ID>
<type>CC_PULSE</type>
<position>-45,-9.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>-25.5,-38.5</position>
<gparam>LABEL_TEXT Accumulator</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-35,-25.5</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>21 </input>
<input>
<ID>IN_2</ID>22 </input>
<input>
<ID>IN_3</ID>23 </input>
<input>
<ID>IN_B_0</ID>19 </input>
<input>
<ID>IN_B_1</ID>19 </input>
<input>
<ID>IN_B_2</ID>19 </input>
<input>
<ID>IN_B_3</ID>19 </input>
<output>
<ID>OUT_0</ID>29 </output>
<output>
<ID>OUT_1</ID>28 </output>
<output>
<ID>OUT_2</ID>27 </output>
<output>
<ID>OUT_3</ID>26 </output>
<input>
<ID>carry_in</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>26</ID>
<type>FF_GND</type>
<position>-4.5,-25.5</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>32</ID>
<type>FF_GND</type>
<position>-25.5,-23</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>38</ID>
<type>AE_REGISTER8</type>
<position>-6,-37</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>32 </input>
<input>
<ID>IN_2</ID>31 </input>
<input>
<ID>IN_3</ID>30 </input>
<input>
<ID>IN_4</ID>29 </input>
<input>
<ID>IN_5</ID>28 </input>
<input>
<ID>IN_6</ID>27 </input>
<input>
<ID>IN_7</ID>26 </input>
<output>
<ID>OUT_0</ID>44 </output>
<output>
<ID>OUT_1</ID>43 </output>
<output>
<ID>OUT_2</ID>42 </output>
<output>
<ID>OUT_3</ID>41 </output>
<output>
<ID>OUT_4</ID>20 </output>
<output>
<ID>OUT_5</ID>21 </output>
<output>
<ID>OUT_6</ID>22 </output>
<output>
<ID>OUT_7</ID>23 </output>
<output>
<ID>carry_out</ID>39 </output>
<input>
<ID>clear</ID>35 </input>
<input>
<ID>clock</ID>34 </input>
<input>
<ID>count_enable</ID>40 </input>
<input>
<ID>count_up</ID>40 </input>
<input>
<ID>load</ID>5 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 97</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>40</ID>
<type>DE_TO</type>
<position>-36.5,-2.5</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>42</ID>
<type>DA_FROM</type>
<position>-9,-43.5</position>
<input>
<ID>IN_0</ID>34 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>44</ID>
<type>DA_FROM</type>
<position>-9,-45.5</position>
<input>
<ID>IN_0</ID>35 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Reset</lparam></gate>
<gate>
<ID>48</ID>
<type>GA_LED</type>
<position>-0.5,-30.5</position>
<input>
<ID>N_in0</ID>39 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>FF_GND</type>
<position>1.5,-29.5</position>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>52</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>12,-37</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>43 </input>
<input>
<ID>IN_2</ID>42 </input>
<input>
<ID>IN_3</ID>41 </input>
<input>
<ID>IN_4</ID>20 </input>
<input>
<ID>IN_5</ID>21 </input>
<input>
<ID>IN_6</ID>22 </input>
<input>
<ID>IN_7</ID>23 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 97</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-18,-1.5,-16.5,-1.5</points>
<connection>
<GID>6</GID>
<name>OUT_2</name></connection>
<connection>
<GID>4</GID>
<name>ADDRESS_2</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-18,-3.5,-16.5,-3.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<connection>
<GID>4</GID>
<name>ADDRESS_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-18,-0.5,-16.5,-0.5</points>
<connection>
<GID>6</GID>
<name>OUT_3</name></connection>
<connection>
<GID>4</GID>
<name>ADDRESS_3</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-18,-2.5,-16.5,-2.5</points>
<connection>
<GID>6</GID>
<name>OUT_1</name></connection>
<connection>
<GID>4</GID>
<name>ADDRESS_1</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-19.5,-31,-7,-31</points>
<connection>
<GID>38</GID>
<name>load</name></connection>
<connection>
<GID>5</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-43,-9.5,-39.5,-9.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5.5,-2.5,-5.5,-1.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6.5,-2.5,-5.5,-2.5</points>
<connection>
<GID>4</GID>
<name>ENABLE_0</name></connection>
<intersection>-5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,5.5,-23,7.5</points>
<connection>
<GID>6</GID>
<name>load</name></connection>
<intersection>7.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-24.5,7.5,-23,7.5</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>-23 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-21,-9,-21,-5.5</points>
<connection>
<GID>6</GID>
<name>clear</name></connection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-21.5,-9,-21,-9</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>-21 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,0.5,-16.5,4</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-18,0.5,-16.5,0.5</points>
<connection>
<GID>6</GID>
<name>OUT_4</name></connection>
<intersection>-16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22,5.5,-22,8</points>
<connection>
<GID>6</GID>
<name>count_enable</name></connection>
<intersection>5.5 3</intersection>
<intersection>8 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-22,8,-13.5,8</points>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-22 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-22,5.5,-21,5.5</points>
<connection>
<GID>6</GID>
<name>count_up</name></connection>
<intersection>-22 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-38.5,-6,-23,-6</points>
<intersection>-38.5 5</intersection>
<intersection>-23 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-23,-6,-23,-5.5</points>
<connection>
<GID>6</GID>
<name>clock</name></connection>
<intersection>-6 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-38.5,-6,-38.5,-2.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>-6 1</intersection>
<intersection>-2.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>-40,-2.5,-38.5,-2.5</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>-38.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27,-24.5,-23,-24.5</points>
<connection>
<GID>24</GID>
<name>carry_in</name></connection>
<connection>
<GID>14</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-21.5,-12,-7</points>
<connection>
<GID>14</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>4</GID>
<name>DATA_OUT_2</name></connection>
<intersection>-10.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-12,-10.5,-9,-10.5</points>
<connection>
<GID>10</GID>
<name>IN_2</name></connection>
<intersection>-12 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,-21.5,-11,-7</points>
<connection>
<GID>14</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>4</GID>
<name>DATA_OUT_1</name></connection>
<intersection>-11.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-11,-11.5,-9,-11.5</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>-11 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13,-21.5,-13,-7</points>
<connection>
<GID>14</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>4</GID>
<name>DATA_OUT_3</name></connection>
<intersection>-9.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-13,-9.5,-9,-9.5</points>
<connection>
<GID>10</GID>
<name>IN_3</name></connection>
<intersection>-13 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,-21.5,-10,-7</points>
<connection>
<GID>14</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>4</GID>
<name>DATA_OUT_0</name></connection>
<intersection>-12.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-10,-12.5,-9,-12.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>-10 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-7,-24.5,-4.5,-24.5</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<connection>
<GID>14</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25.5,-22,-25.5,-21.5</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-33,-21.5,-25.5,-21.5</points>
<connection>
<GID>24</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>24</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>24</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>24</GID>
<name>IN_B_0</name></connection>
<intersection>-25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-21.5,-37,-16.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-37,-16.5,4.5,-16.5</points>
<intersection>-37 0</intersection>
<intersection>4.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>4.5,-36,4.5,-16.5</points>
<intersection>-36 3</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-2,-36,7,-36</points>
<connection>
<GID>38</GID>
<name>OUT_4</name></connection>
<connection>
<GID>52</GID>
<name>IN_4</name></connection>
<intersection>4.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-38,-21.5,-38,-16</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-38,-16,5,-16</points>
<intersection>-38 0</intersection>
<intersection>5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>5,-35,5,-16</points>
<intersection>-35 3</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-2,-35,7,-35</points>
<connection>
<GID>38</GID>
<name>OUT_5</name></connection>
<connection>
<GID>52</GID>
<name>IN_5</name></connection>
<intersection>5 2</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-39,-21.5,-39,-15.5</points>
<connection>
<GID>24</GID>
<name>IN_2</name></connection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-39,-15.5,5.5,-15.5</points>
<intersection>-39 0</intersection>
<intersection>5.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>5.5,-34,5.5,-15.5</points>
<intersection>-34 3</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-2,-34,7,-34</points>
<connection>
<GID>38</GID>
<name>OUT_6</name></connection>
<connection>
<GID>52</GID>
<name>IN_6</name></connection>
<intersection>5.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40,-21.5,-40,-15</points>
<connection>
<GID>24</GID>
<name>IN_3</name></connection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-40,-15,6.5,-15</points>
<intersection>-40 0</intersection>
<intersection>6.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>6.5,-33,6.5,-15</points>
<intersection>-33 3</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-2,-33,7,-33</points>
<connection>
<GID>38</GID>
<name>OUT_7</name></connection>
<connection>
<GID>52</GID>
<name>IN_7</name></connection>
<intersection>6.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,-33,-36.5,-29.5</points>
<connection>
<GID>24</GID>
<name>OUT_3</name></connection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36.5,-33,-10,-33</points>
<connection>
<GID>38</GID>
<name>IN_7</name></connection>
<intersection>-36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-34,-35.5,-29.5</points>
<connection>
<GID>24</GID>
<name>OUT_2</name></connection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35.5,-34,-10,-34</points>
<connection>
<GID>38</GID>
<name>IN_6</name></connection>
<intersection>-35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34.5,-35,-34.5,-29.5</points>
<connection>
<GID>24</GID>
<name>OUT_1</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34.5,-35,-10,-35</points>
<connection>
<GID>38</GID>
<name>IN_5</name></connection>
<intersection>-34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33.5,-36,-33.5,-29.5</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-33.5,-36,-10,-36</points>
<connection>
<GID>38</GID>
<name>IN_4</name></connection>
<intersection>-33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-37,-16.5,-29.5</points>
<connection>
<GID>14</GID>
<name>OUT_3</name></connection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16.5,-37,-10,-37</points>
<connection>
<GID>38</GID>
<name>IN_3</name></connection>
<intersection>-16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15.5,-38,-15.5,-29.5</points>
<connection>
<GID>14</GID>
<name>OUT_2</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15.5,-38,-10,-38</points>
<connection>
<GID>38</GID>
<name>IN_2</name></connection>
<intersection>-15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-39,-14.5,-29.5</points>
<connection>
<GID>14</GID>
<name>OUT_1</name></connection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,-39,-10,-39</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,-40,-13.5,-29.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13.5,-40,-10,-40</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>-13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7,-43.5,-7,-42</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<connection>
<GID>38</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-45.5,-5,-42</points>
<connection>
<GID>38</GID>
<name>clear</name></connection>
<intersection>-45.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7,-45.5,-5,-45.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>-5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-31,-4,-30.5</points>
<connection>
<GID>38</GID>
<name>carry_out</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4,-30.5,-1.5,-30.5</points>
<connection>
<GID>48</GID>
<name>N_in0</name></connection>
<intersection>-4 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-31,-5,-28.5</points>
<connection>
<GID>38</GID>
<name>count_up</name></connection>
<intersection>-31 4</intersection>
<intersection>-28.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-5,-28.5,1.5,-28.5</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>-5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-6,-31,-5,-31</points>
<connection>
<GID>38</GID>
<name>count_enable</name></connection>
<intersection>-5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-37,7,-37</points>
<connection>
<GID>38</GID>
<name>OUT_3</name></connection>
<connection>
<GID>52</GID>
<name>IN_3</name></connection>
<intersection>4 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>4,-37,4,-17</points>
<intersection>-37 1</intersection>
<intersection>-17 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-20,-17,4,-17</points>
<intersection>-20 9</intersection>
<intersection>4 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-20,-21.5,-20,-17</points>
<connection>
<GID>14</GID>
<name>IN_3</name></connection>
<intersection>-17 8</intersection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-38,7,-38</points>
<connection>
<GID>38</GID>
<name>OUT_2</name></connection>
<connection>
<GID>52</GID>
<name>IN_2</name></connection>
<intersection>3.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>3.5,-38,3.5,-17.5</points>
<intersection>-38 1</intersection>
<intersection>-17.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-19,-17.5,3.5,-17.5</points>
<intersection>-19 9</intersection>
<intersection>3.5 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-19,-21.5,-19,-17.5</points>
<connection>
<GID>14</GID>
<name>IN_2</name></connection>
<intersection>-17.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-39,7,-39</points>
<connection>
<GID>38</GID>
<name>OUT_1</name></connection>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>3 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>3,-39,3,-18</points>
<intersection>-39 1</intersection>
<intersection>-18 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-18,-18,3,-18</points>
<intersection>-18 9</intersection>
<intersection>3 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-18,-21.5,-18,-18</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>-18 8</intersection></vsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-40,7,-40</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>2.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>2.5,-40,2.5,-18.5</points>
<intersection>-40 1</intersection>
<intersection>-18.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-17,-18.5,2.5,-18.5</points>
<intersection>-17 9</intersection>
<intersection>2.5 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-17,-21.5,-17,-18.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>-18.5 8</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>13.5705,21.3384,189.903,-100.215</PageViewport></page 1>
<page 2>
<PageViewport>-5.37044,44.0087,314.324,-176.37</PageViewport></page 2>
<page 3>
<PageViewport>-5.37044,44.0087,314.324,-176.37</PageViewport></page 3>
<page 4>
<PageViewport>-5.37044,44.0087,314.324,-176.37</PageViewport></page 4>
<page 5>
<PageViewport>-5.37044,44.0087,314.324,-176.37</PageViewport></page 5>
<page 6>
<PageViewport>-5.37044,44.0087,314.324,-176.37</PageViewport></page 6>
<page 7>
<PageViewport>-5.37044,44.0087,314.324,-176.37</PageViewport></page 7>
<page 8>
<PageViewport>-5.37044,44.0087,314.324,-176.37</PageViewport></page 8>
<page 9>
<PageViewport>-5.37044,44.0087,314.324,-176.37</PageViewport></page 9></circuit>