<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-5.02458,50.938,110.449,-15.25</PageViewport>
<gate>
<ID>2</ID>
<type>DE_TO</type>
<position>7.5,44.5</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>81,48</position>
<gparam>LABEL_TEXT Alex Laird</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>DE_TO</type>
<position>7.5,41.5</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_LABEL</type>
<position>81,44.5</position>
<gparam>LABEL_TEXT Gates Used: 14</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>DE_TO</type>
<position>7.5,38.5</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>81,41</position>
<gparam>LABEL_TEXT Inputs: 41</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>DE_TO</type>
<position>7.5,35.5</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>81,37.5</position>
<gparam>LABEL_TEXT Cost = 83</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>3.5,44.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_TOGGLE</type>
<position>3.5,41.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>3.5,38.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_TOGGLE</type>
<position>3.5,35.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>15</ID>
<type>DA_FROM</type>
<position>15,44.5</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>16</ID>
<type>DA_FROM</type>
<position>15,42.5</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>18</ID>
<type>DA_FROM</type>
<position>15,40</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>19</ID>
<type>DA_FROM</type>
<position>15,38</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>20</ID>
<type>DA_FROM</type>
<position>15,36</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>21</ID>
<type>DA_FROM</type>
<position>15,33.5</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>22</ID>
<type>DA_FROM</type>
<position>15,31.5</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>23</ID>
<type>DA_FROM</type>
<position>15,29.5</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>25</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,38</position>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,33.5</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>27</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,31.5</position>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>28</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,29.5</position>
<input>
<ID>IN_0</ID>8 </input>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_AND3</type>
<position>24,38</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>9 </input>
<input>
<ID>IN_2</ID>14 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_AND3</type>
<position>24,31.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<input>
<ID>IN_2</ID>12 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>34</ID>
<type>AE_OR4</type>
<position>34.5,41.5</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>16 </input>
<input>
<ID>IN_2</ID>17 </input>
<input>
<ID>IN_3</ID>18 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>35</ID>
<type>DE_TO</type>
<position>42.5,41.5</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID a</lparam></gate>
<gate>
<ID>36</ID>
<type>DE_TO</type>
<position>35.5,34.5</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BC'D</lparam></gate>
<gate>
<ID>37</ID>
<type>DE_TO</type>
<position>35.5,32.5</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B'C'D'</lparam></gate>
<gate>
<ID>38</ID>
<type>DA_FROM</type>
<position>15,25.5</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>39</ID>
<type>DA_FROM</type>
<position>15,23.5</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>40</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,23.5</position>
<input>
<ID>IN_0</ID>20 </input>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>42</ID>
<type>AO_XNOR2</type>
<position>20,20</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>22 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>43</ID>
<type>DA_FROM</type>
<position>15,21</position>
<input>
<ID>IN_0</ID>21 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>44</ID>
<type>DA_FROM</type>
<position>15,19</position>
<input>
<ID>IN_0</ID>22 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>46</ID>
<type>AE_OR3</type>
<position>28,23.5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>25 </input>
<input>
<ID>IN_2</ID>23 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>47</ID>
<type>DE_TO</type>
<position>35,23.5</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID b</lparam></gate>
<gate>
<ID>48</ID>
<type>DA_FROM</type>
<position>15,15</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>49</ID>
<type>DA_FROM</type>
<position>15,13</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>50</ID>
<type>DA_FROM</type>
<position>15,11</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>51</ID>
<type>DA_FROM</type>
<position>15,9</position>
<input>
<ID>IN_0</ID>31 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>53</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,11</position>
<input>
<ID>IN_0</ID>27 </input>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>54</ID>
<type>AE_OR4</type>
<position>24,12</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>30 </input>
<input>
<ID>IN_2</ID>28 </input>
<input>
<ID>IN_3</ID>31 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>55</ID>
<type>DE_TO</type>
<position>32,12</position>
<input>
<ID>IN_0</ID>32 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID c</lparam></gate>
<gate>
<ID>56</ID>
<type>DA_FROM</type>
<position>15,5</position>
<input>
<ID>IN_0</ID>39 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>57</ID>
<type>DA_FROM</type>
<position>15,3</position>
<input>
<ID>IN_0</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B'C'D'</lparam></gate>
<gate>
<ID>58</ID>
<type>DA_FROM</type>
<position>15,-1.5</position>
<input>
<ID>IN_0</ID>35 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>59</ID>
<type>DA_FROM</type>
<position>15,-3.5</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>60</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,-3.5</position>
<input>
<ID>IN_0</ID>33 </input>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_AND2</type>
<position>24,-2.5</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>63</ID>
<type>DA_FROM</type>
<position>15,-6</position>
<input>
<ID>IN_0</ID>36 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>64</ID>
<type>DA_FROM</type>
<position>15,-8</position>
<input>
<ID>IN_0</ID>38 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>65</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,-6</position>
<input>
<ID>IN_0</ID>36 </input>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_AND2</type>
<position>24,-7</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>67</ID>
<type>DA_FROM</type>
<position>15,1</position>
<input>
<ID>IN_0</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BC'D</lparam></gate>
<gate>
<ID>69</ID>
<type>DE_OR8</type>
<position>34.5,1.5</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>40 </input>
<input>
<ID>IN_2</ID>41 </input>
<input>
<ID>IN_3</ID>42 </input>
<input>
<ID>IN_4</ID>43 </input>
<input>
<ID>IN_5</ID>43 </input>
<input>
<ID>IN_6</ID>43 </input>
<input>
<ID>IN_7</ID>43 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>70</ID>
<type>DE_TO</type>
<position>34,-5.5</position>
<input>
<ID>IN_0</ID>42 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CD'</lparam></gate>
<gate>
<ID>71</ID>
<type>DE_TO</type>
<position>40.5,1.5</position>
<input>
<ID>IN_0</ID>44 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID d</lparam></gate>
<gate>
<ID>72</ID>
<type>DA_FROM</type>
<position>15,-12</position>
<input>
<ID>IN_0</ID>45 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CD'</lparam></gate>
<gate>
<ID>73</ID>
<type>DA_FROM</type>
<position>15,-14</position>
<input>
<ID>IN_0</ID>46 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B'C'D'</lparam></gate>
<gate>
<ID>75</ID>
<type>AE_OR2</type>
<position>21.5,-13</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>DE_TO</type>
<position>28,-13</position>
<input>
<ID>IN_0</ID>47 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID e</lparam></gate>
<gate>
<ID>77</ID>
<type>DA_FROM</type>
<position>47,19.5</position>
<input>
<ID>IN_0</ID>55 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>78</ID>
<type>DA_FROM</type>
<position>47,17.5</position>
<input>
<ID>IN_0</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BC'D</lparam></gate>
<gate>
<ID>79</ID>
<type>DA_FROM</type>
<position>47,15</position>
<input>
<ID>IN_0</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>80</ID>
<type>DA_FROM</type>
<position>47,13</position>
<input>
<ID>IN_0</ID>50 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>81</ID>
<type>DA_FROM</type>
<position>47,10.5</position>
<input>
<ID>IN_0</ID>54 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>82</ID>
<type>DA_FROM</type>
<position>47,8.5</position>
<input>
<ID>IN_0</ID>48 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>83</ID>
<type>AE_SMALL_INVERTER</type>
<position>51,8.5</position>
<input>
<ID>IN_0</ID>48 </input>
<output>
<ID>OUT_0</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>84</ID>
<type>AE_SMALL_INVERTER</type>
<position>51,15</position>
<input>
<ID>IN_0</ID>49 </input>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>85</ID>
<type>AE_SMALL_INVERTER</type>
<position>51,13</position>
<input>
<ID>IN_0</ID>50 </input>
<output>
<ID>OUT_0</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>87</ID>
<type>AA_AND2</type>
<position>56,14</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>52 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>89</ID>
<type>AA_AND2</type>
<position>56,9.5</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>53 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>91</ID>
<type>AE_OR4</type>
<position>65,16.5</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>56 </input>
<input>
<ID>IN_2</ID>57 </input>
<input>
<ID>IN_3</ID>58 </input>
<output>
<ID>OUT</ID>59 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>92</ID>
<type>DE_TO</type>
<position>72.5,16.5</position>
<input>
<ID>IN_0</ID>59 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID f</lparam></gate>
<gate>
<ID>93</ID>
<type>DA_FROM</type>
<position>47,4.5</position>
<input>
<ID>IN_0</ID>60 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>94</ID>
<type>DA_FROM</type>
<position>47,2.5</position>
<input>
<ID>IN_0</ID>61 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>95</ID>
<type>DA_FROM</type>
<position>47,0.5</position>
<input>
<ID>IN_0</ID>62 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>97</ID>
<type>AE_OR3</type>
<position>53.5,2.5</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>61 </input>
<input>
<ID>IN_2</ID>62 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>98</ID>
<type>DE_TO</type>
<position>60,2.5</position>
<input>
<ID>IN_0</ID>63 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID g</lparam></gate>
<gate>
<ID>100</ID>
<type>GA_LED</type>
<position>52.5,44.5</position>
<input>
<ID>N_in2</ID>64 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>101</ID>
<type>GA_LED</type>
<position>52.5,42.5</position>
<input>
<ID>N_in0</ID>93 </input>
<input>
<ID>N_in2</ID>65 </input>
<input>
<ID>N_in3</ID>64 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>102</ID>
<type>GA_LED</type>
<position>52.5,40.5</position>
<input>
<ID>N_in2</ID>66 </input>
<input>
<ID>N_in3</ID>65 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>103</ID>
<type>GA_LED</type>
<position>52.5,38.5</position>
<input>
<ID>N_in3</ID>66 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>104</ID>
<type>GA_LED</type>
<position>54.5,46.5</position>
<input>
<ID>N_in1</ID>67 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>GA_LED</type>
<position>56.5,46.5</position>
<input>
<ID>N_in0</ID>67 </input>
<input>
<ID>N_in1</ID>68 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>106</ID>
<type>GA_LED</type>
<position>58.5,46.5</position>
<input>
<ID>N_in0</ID>68 </input>
<input>
<ID>N_in1</ID>69 </input>
<input>
<ID>N_in3</ID>88 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>107</ID>
<type>GA_LED</type>
<position>60.5,46.5</position>
<input>
<ID>N_in0</ID>69 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>GA_LED</type>
<position>62.5,44.5</position>
<input>
<ID>N_in2</ID>70 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>109</ID>
<type>GA_LED</type>
<position>62.5,42.5</position>
<input>
<ID>N_in1</ID>89 </input>
<input>
<ID>N_in2</ID>71 </input>
<input>
<ID>N_in3</ID>70 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>GA_LED</type>
<position>62.5,40.5</position>
<input>
<ID>N_in2</ID>72 </input>
<input>
<ID>N_in3</ID>71 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>GA_LED</type>
<position>62.5,38.5</position>
<input>
<ID>N_in3</ID>72 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>112</ID>
<type>GA_LED</type>
<position>60.5,36.5</position>
<input>
<ID>N_in0</ID>73 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>113</ID>
<type>GA_LED</type>
<position>58.5,36.5</position>
<input>
<ID>N_in0</ID>74 </input>
<input>
<ID>N_in1</ID>73 </input>
<input>
<ID>N_in3</ID>87 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>GA_LED</type>
<position>56.5,36.5</position>
<input>
<ID>N_in0</ID>86 </input>
<input>
<ID>N_in1</ID>74 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>115</ID>
<type>GA_LED</type>
<position>54.5,36.5</position>
<input>
<ID>N_in1</ID>86 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>GA_LED</type>
<position>52.5,34.5</position>
<input>
<ID>N_in2</ID>76 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>GA_LED</type>
<position>52.5,32.5</position>
<input>
<ID>N_in0</ID>92 </input>
<input>
<ID>N_in2</ID>77 </input>
<input>
<ID>N_in3</ID>76 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>119</ID>
<type>GA_LED</type>
<position>52.5,30.5</position>
<input>
<ID>N_in2</ID>82 </input>
<input>
<ID>N_in3</ID>77 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>120</ID>
<type>GA_LED</type>
<position>62.5,34.5</position>
<input>
<ID>N_in2</ID>78 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>121</ID>
<type>GA_LED</type>
<position>62.5,32.5</position>
<input>
<ID>N_in1</ID>90 </input>
<input>
<ID>N_in2</ID>79 </input>
<input>
<ID>N_in3</ID>78 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>GA_LED</type>
<position>62.5,30.5</position>
<input>
<ID>N_in2</ID>80 </input>
<input>
<ID>N_in3</ID>79 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>123</ID>
<type>GA_LED</type>
<position>62.5,28.5</position>
<input>
<ID>N_in3</ID>80 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>125</ID>
<type>GA_LED</type>
<position>52.5,28.5</position>
<input>
<ID>N_in3</ID>82 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>126</ID>
<type>GA_LED</type>
<position>54.5,26.5</position>
<input>
<ID>N_in1</ID>83 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>127</ID>
<type>GA_LED</type>
<position>56.5,26.5</position>
<input>
<ID>N_in0</ID>83 </input>
<input>
<ID>N_in1</ID>84 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>GA_LED</type>
<position>58.5,26.5</position>
<input>
<ID>N_in0</ID>84 </input>
<input>
<ID>N_in1</ID>85 </input>
<input>
<ID>N_in2</ID>91 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>GA_LED</type>
<position>60.5,26.5</position>
<input>
<ID>N_in0</ID>85 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>DA_FROM</type>
<position>58.5,39.5</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID g</lparam></gate>
<gate>
<ID>131</ID>
<type>DA_FROM</type>
<position>58.5,49.5</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID a</lparam></gate>
<gate>
<ID>132</ID>
<type>DA_FROM</type>
<position>65.5,42.5</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID b</lparam></gate>
<gate>
<ID>133</ID>
<type>DA_FROM</type>
<position>65.5,32.5</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID c</lparam></gate>
<gate>
<ID>134</ID>
<type>DA_FROM</type>
<position>58.5,23.5</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID d</lparam></gate>
<gate>
<ID>135</ID>
<type>DA_FROM</type>
<position>49.5,32.5</position>
<input>
<ID>IN_0</ID>92 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID e</lparam></gate>
<gate>
<ID>136</ID>
<type>DA_FROM</type>
<position>49.5,42.5</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID f</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,44.5,5.5,44.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,41.5,5.5,41.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,38.5,5.5,38.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,35.5,5.5,35.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,38,17,38</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<connection>
<GID>25</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,33.5,17,33.5</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<connection>
<GID>26</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,31.5,17,31.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<connection>
<GID>27</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,29.5,17,29.5</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<connection>
<GID>28</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,38,21,38</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<connection>
<GID>30</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,33.5,21,33.5</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<connection>
<GID>32</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,31.5,21,31.5</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<connection>
<GID>32</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,29.5,21,29.5</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<connection>
<GID>32</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,40,21,40</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<connection>
<GID>18</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,36,21,36</points>
<connection>
<GID>30</GID>
<name>IN_2</name></connection>
<connection>
<GID>20</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,44.5,31.5,44.5</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<connection>
<GID>34</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,42.5,31.5,42.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<connection>
<GID>34</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,34.5,29,40.5</points>
<intersection>34.5 3</intersection>
<intersection>38 2</intersection>
<intersection>40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,40.5,31.5,40.5</points>
<connection>
<GID>34</GID>
<name>IN_2</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,38,29,38</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>29,34.5,33.5,34.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,31.5,30,38.5</points>
<intersection>31.5 2</intersection>
<intersection>32.5 3</intersection>
<intersection>38.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,38.5,31.5,38.5</points>
<connection>
<GID>34</GID>
<name>IN_3</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,31.5,30,31.5</points>
<connection>
<GID>32</GID>
<name>OUT</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30,32.5,33.5,32.5</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38.5,41.5,40.5,41.5</points>
<connection>
<GID>34</GID>
<name>OUT</name></connection>
<connection>
<GID>35</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,23.5,17,23.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<connection>
<GID>40</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,21,17,21</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<connection>
<GID>43</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,19,17,19</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<connection>
<GID>44</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,21.5,25,21.5</points>
<connection>
<GID>46</GID>
<name>IN_2</name></connection>
<intersection>24 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>24,20,24,21.5</points>
<intersection>20 5</intersection>
<intersection>21.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>23,20,24,20</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<intersection>24 4</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,25.5,25,25.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<connection>
<GID>46</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21,23.5,25,23.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<connection>
<GID>46</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,23.5,33,23.5</points>
<connection>
<GID>46</GID>
<name>OUT</name></connection>
<connection>
<GID>47</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,11,17,11</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<connection>
<GID>53</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,11,21,11</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<connection>
<GID>54</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,15,21,15</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<connection>
<GID>48</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,13,21,13</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<connection>
<GID>49</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,9,21,9</points>
<connection>
<GID>54</GID>
<name>IN_3</name></connection>
<connection>
<GID>51</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28,12,30,12</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<connection>
<GID>55</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-3.5,17,-3.5</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<connection>
<GID>60</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-3.5,21,-3.5</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<connection>
<GID>62</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,-1.5,21,-1.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<connection>
<GID>58</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-6,17,-6</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<connection>
<GID>65</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-6,21,-6</points>
<connection>
<GID>65</GID>
<name>OUT_0</name></connection>
<connection>
<GID>66</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,-8,21,-8</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<connection>
<GID>64</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,5,31.5,5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<connection>
<GID>56</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,3,24,4</points>
<intersection>3 2</intersection>
<intersection>4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,4,31.5,4</points>
<connection>
<GID>69</GID>
<name>IN_1</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,3,24,3</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,1,25,3</points>
<intersection>1 2</intersection>
<intersection>3 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,3,31.5,3</points>
<connection>
<GID>69</GID>
<name>IN_2</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,1,25,1</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-5.5,28,2</points>
<intersection>-5.5 3</intersection>
<intersection>-2.5 2</intersection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,2,31.5,2</points>
<connection>
<GID>69</GID>
<name>IN_3</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-2.5,28,-2.5</points>
<connection>
<GID>62</GID>
<name>OUT</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>28,-5.5,32,-5.5</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-7,29,1</points>
<intersection>-7 2</intersection>
<intersection>1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,1,31.5,1</points>
<connection>
<GID>69</GID>
<name>IN_7</name></connection>
<intersection>29 0</intersection>
<intersection>31.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-7,29,-7</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<intersection>29 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>31.5,-2,31.5,1</points>
<connection>
<GID>69</GID>
<name>IN_4</name></connection>
<connection>
<GID>69</GID>
<name>IN_6</name></connection>
<connection>
<GID>69</GID>
<name>IN_5</name></connection>
<intersection>1 1</intersection></vsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,1.5,38.5,1.5</points>
<connection>
<GID>69</GID>
<name>OUT</name></connection>
<connection>
<GID>71</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,-12,18.5,-12</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<connection>
<GID>75</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,-14,18.5,-14</points>
<connection>
<GID>75</GID>
<name>IN_1</name></connection>
<connection>
<GID>73</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-13,26,-13</points>
<connection>
<GID>75</GID>
<name>OUT</name></connection>
<connection>
<GID>76</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,8.5,49,8.5</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<connection>
<GID>83</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,15,49,15</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<connection>
<GID>84</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,13,49,13</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<connection>
<GID>85</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,15,53,15</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<connection>
<GID>87</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,13,53,13</points>
<connection>
<GID>85</GID>
<name>OUT_0</name></connection>
<connection>
<GID>87</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,8.5,53,8.5</points>
<connection>
<GID>83</GID>
<name>OUT_0</name></connection>
<connection>
<GID>89</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49,10.5,53,10.5</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<connection>
<GID>81</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49,19.5,62,19.5</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<connection>
<GID>77</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49,17.5,62,17.5</points>
<connection>
<GID>91</GID>
<name>IN_1</name></connection>
<connection>
<GID>78</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,14,60,15.5</points>
<intersection>14 2</intersection>
<intersection>15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60,15.5,62,15.5</points>
<connection>
<GID>91</GID>
<name>IN_2</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59,14,60,14</points>
<connection>
<GID>87</GID>
<name>OUT</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,9.5,61,13.5</points>
<intersection>9.5 2</intersection>
<intersection>13.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>59,9.5,61,9.5</points>
<connection>
<GID>89</GID>
<name>OUT</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>61,13.5,62,13.5</points>
<connection>
<GID>91</GID>
<name>IN_3</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69,16.5,70.5,16.5</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<connection>
<GID>91</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49,4.5,50.5,4.5</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<connection>
<GID>93</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49,2.5,50.5,2.5</points>
<connection>
<GID>97</GID>
<name>IN_1</name></connection>
<connection>
<GID>94</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49,0.5,50.5,0.5</points>
<connection>
<GID>97</GID>
<name>IN_2</name></connection>
<connection>
<GID>95</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56.5,2.5,58,2.5</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<connection>
<GID>97</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,43.5,52.5,43.5</points>
<connection>
<GID>100</GID>
<name>N_in2</name></connection>
<connection>
<GID>101</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,41.5,52.5,41.5</points>
<connection>
<GID>101</GID>
<name>N_in2</name></connection>
<connection>
<GID>102</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,39.5,52.5,39.5</points>
<connection>
<GID>102</GID>
<name>N_in2</name></connection>
<connection>
<GID>103</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,46.5,55.5,46.5</points>
<connection>
<GID>104</GID>
<name>N_in1</name></connection>
<connection>
<GID>105</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,46.5,57.5,46.5</points>
<connection>
<GID>105</GID>
<name>N_in1</name></connection>
<connection>
<GID>106</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,46.5,59.5,46.5</points>
<connection>
<GID>106</GID>
<name>N_in1</name></connection>
<connection>
<GID>107</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,43.5,62.5,43.5</points>
<connection>
<GID>108</GID>
<name>N_in2</name></connection>
<connection>
<GID>109</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,41.5,62.5,41.5</points>
<connection>
<GID>109</GID>
<name>N_in2</name></connection>
<connection>
<GID>110</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,39.5,62.5,39.5</points>
<connection>
<GID>110</GID>
<name>N_in2</name></connection>
<connection>
<GID>111</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,36.5,59.5,36.5</points>
<connection>
<GID>112</GID>
<name>N_in0</name></connection>
<connection>
<GID>113</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,36.5,57.5,36.5</points>
<connection>
<GID>113</GID>
<name>N_in0</name></connection>
<connection>
<GID>114</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,33.5,52.5,33.5</points>
<connection>
<GID>116</GID>
<name>N_in2</name></connection>
<connection>
<GID>118</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,31.5,52.5,31.5</points>
<connection>
<GID>118</GID>
<name>N_in2</name></connection>
<connection>
<GID>119</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,33.5,62.5,33.5</points>
<connection>
<GID>120</GID>
<name>N_in2</name></connection>
<connection>
<GID>121</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,31.5,62.5,31.5</points>
<connection>
<GID>121</GID>
<name>N_in2</name></connection>
<connection>
<GID>122</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,29.5,62.5,29.5</points>
<connection>
<GID>122</GID>
<name>N_in2</name></connection>
<connection>
<GID>123</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,29.5,52.5,29.5</points>
<connection>
<GID>119</GID>
<name>N_in2</name></connection>
<connection>
<GID>125</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,26.5,55.5,26.5</points>
<connection>
<GID>126</GID>
<name>N_in1</name></connection>
<connection>
<GID>127</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,26.5,57.5,26.5</points>
<connection>
<GID>127</GID>
<name>N_in1</name></connection>
<connection>
<GID>128</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,26.5,59.5,26.5</points>
<connection>
<GID>128</GID>
<name>N_in1</name></connection>
<connection>
<GID>129</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,36.5,55.5,36.5</points>
<connection>
<GID>114</GID>
<name>N_in0</name></connection>
<connection>
<GID>115</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,37.5,58.5,37.5</points>
<connection>
<GID>113</GID>
<name>N_in3</name></connection>
<connection>
<GID>130</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,47.5,58.5,47.5</points>
<connection>
<GID>106</GID>
<name>N_in3</name></connection>
<connection>
<GID>131</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,42.5,63.5,42.5</points>
<connection>
<GID>109</GID>
<name>N_in1</name></connection>
<connection>
<GID>132</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,32.5,63.5,32.5</points>
<connection>
<GID>121</GID>
<name>N_in1</name></connection>
<connection>
<GID>133</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,25.5,58.5,25.5</points>
<connection>
<GID>128</GID>
<name>N_in2</name></connection>
<connection>
<GID>134</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,32.5,51.5,32.5</points>
<connection>
<GID>118</GID>
<name>N_in0</name></connection>
<connection>
<GID>135</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,42.5,51.5,42.5</points>
<connection>
<GID>101</GID>
<name>N_in0</name></connection>
<connection>
<GID>136</GID>
<name>IN_0</name></connection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>-1.24625,31.151,380.343,-187.572</PageViewport></page 1>
<page 2>
<PageViewport>-1.24625,31.151,380.343,-187.572</PageViewport></page 2>
<page 3>
<PageViewport>-1.24625,31.151,380.343,-187.572</PageViewport></page 3>
<page 4>
<PageViewport>-1.24625,31.151,380.343,-187.572</PageViewport></page 4>
<page 5>
<PageViewport>-1.24625,31.151,380.343,-187.572</PageViewport></page 5>
<page 6>
<PageViewport>-1.24625,31.151,380.343,-187.572</PageViewport></page 6>
<page 7>
<PageViewport>-1.24625,31.151,380.343,-187.572</PageViewport></page 7>
<page 8>
<PageViewport>-1.24625,31.151,380.343,-187.572</PageViewport></page 8>
<page 9>
<PageViewport>-1.24625,31.151,380.343,-187.572</PageViewport></page 9></circuit>