<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>14.6642,-13.269,85.2545,-62.25</PageViewport>
<gate>
<ID>2</ID>
<type>DD_KEYPAD_HEX</type>
<position>23.5,-23</position>
<output>
<ID>OUT_0</ID>4 </output>
<output>
<ID>OUT_1</ID>3 </output>
<output>
<ID>OUT_2</ID>2 </output>
<output>
<ID>OUT_3</ID>1 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 14</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>57.5,-31</position>
<gparam>LABEL_TEXT Subtract/Add</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>38,-23</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>2 </input>
<input>
<ID>IN_3</ID>1 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 14</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>6</ID>
<type>AE_FULLADDER_4BIT</type>
<position>35,-51</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>2 </input>
<input>
<ID>IN_3</ID>1 </input>
<input>
<ID>IN_B_0</ID>13 </input>
<input>
<ID>IN_B_1</ID>12 </input>
<input>
<ID>IN_B_2</ID>11 </input>
<input>
<ID>IN_B_3</ID>10 </input>
<output>
<ID>OUT_0</ID>23 </output>
<output>
<ID>OUT_1</ID>22 </output>
<output>
<ID>OUT_2</ID>21 </output>
<output>
<ID>OUT_3</ID>20 </output>
<input>
<ID>carry_in</ID>18 </input>
<output>
<ID>overflow</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>7</ID>
<type>DD_KEYPAD_HEX</type>
<position>45,-23</position>
<output>
<ID>OUT_0</ID>17 </output>
<output>
<ID>OUT_1</ID>16 </output>
<output>
<ID>OUT_2</ID>15 </output>
<output>
<ID>OUT_3</ID>14 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 6</lparam></gate>
<gate>
<ID>8</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>58,-23</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>16 </input>
<input>
<ID>IN_2</ID>15 </input>
<input>
<ID>IN_3</ID>14 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 6</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>47.5,-52.5</position>
<gparam>LABEL_TEXT Note: Numbers >7 are negative</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>48,-54.5</position>
<gparam>LABEL_TEXT 8=-8, 9=-7, A=-6, B=-5</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>48,-56.5</position>
<gparam>LABEL_TEXT C=-4, D=-3, E=-2, F=-1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AI_XOR2</type>
<position>50.5,-38.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>AI_XOR2</type>
<position>46,-38.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AI_XOR2</type>
<position>41.5,-38.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>AI_XOR2</type>
<position>37,-38.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_TOGGLE</type>
<position>64.5,-34</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>20,-14.5</position>
<gparam>LABEL_TEXT 2's Complement Adder Subtracter</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>40.5,-59</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>22 </input>
<input>
<ID>IN_2</ID>21 </input>
<input>
<ID>IN_3</ID>20 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 4</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>18.5,-54</position>
<gparam>LABEL_TEXT Overflow</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>GA_LED</type>
<position>24.5,-52</position>
<input>
<ID>N_in1</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-21,28.5,-20</points>
<connection>
<GID>2</GID>
<name>OUT_3</name></connection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-21,35,-21</points>
<connection>
<GID>4</GID>
<name>IN_3</name></connection>
<intersection>28.5 0</intersection>
<intersection>30 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>30,-47,30,-21</points>
<connection>
<GID>6</GID>
<name>IN_3</name></connection>
<intersection>-21 2</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>28.5,-22,35,-22</points>
<connection>
<GID>2</GID>
<name>OUT_2</name></connection>
<connection>
<GID>4</GID>
<name>IN_2</name></connection>
<intersection>31 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31,-47,31,-22</points>
<connection>
<GID>6</GID>
<name>IN_2</name></connection>
<intersection>-22 2</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-24,28.5,-23</points>
<connection>
<GID>2</GID>
<name>OUT_1</name></connection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-23,35,-23</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>28.5 0</intersection>
<intersection>32 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>32,-47,32,-23</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>-23 2</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-47,33,-24</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>-26 1</intersection>
<intersection>-24 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-26,33,-26</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>33,-24,35,-24</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-47,37,-41.5</points>
<connection>
<GID>6</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>15</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-47,38,-44</points>
<connection>
<GID>6</GID>
<name>IN_B_2</name></connection>
<intersection>-44 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>41.5,-44,41.5,-41.5</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>-44 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>38,-44,41.5,-44</points>
<intersection>38 0</intersection>
<intersection>41.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-47,39,-45</points>
<connection>
<GID>6</GID>
<name>IN_B_1</name></connection>
<intersection>-45 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>46,-45,46,-41.5</points>
<connection>
<GID>13</GID>
<name>OUT</name></connection>
<intersection>-45 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>39,-45,46,-45</points>
<intersection>39 0</intersection>
<intersection>46 1</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-47,50.5,-41.5</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>-47 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>40,-47,50.5,-47</points>
<connection>
<GID>6</GID>
<name>IN_B_0</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-30.5,51,-20</points>
<intersection>-30.5 3</intersection>
<intersection>-21 1</intersection>
<intersection>-20 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-21,55,-21</points>
<connection>
<GID>8</GID>
<name>IN_3</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>36,-30.5,51,-30.5</points>
<intersection>36 4</intersection>
<intersection>51 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>36,-35.5,36,-30.5</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>-30.5 3</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>50,-20,51,-20</points>
<connection>
<GID>7</GID>
<name>OUT_3</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-31.5,52,-22</points>
<intersection>-31.5 4</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-22,55,-22</points>
<connection>
<GID>7</GID>
<name>OUT_2</name></connection>
<connection>
<GID>8</GID>
<name>IN_2</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>40.5,-31.5,52,-31.5</points>
<intersection>40.5 5</intersection>
<intersection>52 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>40.5,-35.5,40.5,-31.5</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>-31.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-32.5,53,-23</points>
<intersection>-32.5 3</intersection>
<intersection>-24 10</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-23,55,-23</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>45,-32.5,53,-32.5</points>
<intersection>45 4</intersection>
<intersection>53 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>45,-35.5,45,-32.5</points>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<intersection>-32.5 3</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>50,-24,53,-24</points>
<connection>
<GID>7</GID>
<name>OUT_1</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-34.5,54,-24</points>
<intersection>-34.5 2</intersection>
<intersection>-26 4</intersection>
<intersection>-24 9</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-34.5,54,-34.5</points>
<intersection>49.5 5</intersection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>50,-26,54,-26</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>54 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>49.5,-35.5,49.5,-34.5</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>54,-24,55,-24</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-34,62.5,-34</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<intersection>38 6</intersection>
<intersection>42.5 11</intersection>
<intersection>47 5</intersection>
<intersection>51.5 4</intersection>
<intersection>56 7</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>51.5,-35.5,51.5,-34</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>-34 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>47,-35.5,47,-34</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>-34 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>38,-35.5,38,-34</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>-34 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>56,-50,56,-34</points>
<intersection>-50 9</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>43,-50,56,-50</points>
<connection>
<GID>6</GID>
<name>carry_in</name></connection>
<intersection>56 7</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>42.5,-35.5,42.5,-34</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>-34 1</intersection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-57,33.5,-55</points>
<connection>
<GID>6</GID>
<name>OUT_3</name></connection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-57,37.5,-57</points>
<connection>
<GID>19</GID>
<name>IN_3</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-58,34.5,-55</points>
<connection>
<GID>6</GID>
<name>OUT_2</name></connection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-58,37.5,-58</points>
<connection>
<GID>19</GID>
<name>IN_2</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-59,35.5,-55</points>
<connection>
<GID>6</GID>
<name>OUT_1</name></connection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-59,37.5,-59</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-60,36.5,-55</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-60,37.5,-60</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-52,27,-52</points>
<connection>
<GID>6</GID>
<name>overflow</name></connection>
<connection>
<GID>21</GID>
<name>N_in1</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-1.41973,1.18513,89.6197,-61.9851</PageViewport></page 1>
<page 2>
<PageViewport>-1.41973,1.18513,89.6197,-61.9851</PageViewport></page 2>
<page 3>
<PageViewport>-1.41973,1.18513,89.6197,-61.9851</PageViewport></page 3>
<page 4>
<PageViewport>-1.41973,1.18513,89.6197,-61.9851</PageViewport></page 4>
<page 5>
<PageViewport>-1.41973,1.18513,89.6197,-61.9851</PageViewport></page 5>
<page 6>
<PageViewport>-1.41973,1.18513,89.6197,-61.9851</PageViewport></page 6>
<page 7>
<PageViewport>-1.41973,1.18513,89.6197,-61.9851</PageViewport></page 7>
<page 8>
<PageViewport>-1.41973,1.18513,89.6197,-61.9851</PageViewport></page 8>
<page 9>
<PageViewport>-1.41973,1.18513,89.6197,-61.9851</PageViewport></page 9></circuit>