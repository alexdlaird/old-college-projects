<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-18.0092,25.25,99.7529,-42.25</PageViewport>
<gate>
<ID>2</ID>
<type>AA_AND3</type>
<position>8.5,-8</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>17 </input>
<input>
<ID>IN_2</ID>18 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>3</ID>
<type>BI_NANDX3</type>
<position>62,-14</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>31 </input>
<input>
<ID>IN_2</ID>30 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_AND2</type>
<position>8.5,-14</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_AND2</type>
<position>8,-19</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>BM_NORX3</type>
<position>60,-35</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>41 </input>
<input>
<ID>IN_2</ID>42 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>7</ID>
<type>AE_OR3</type>
<position>22,-14</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>4 </input>
<input>
<ID>IN_2</ID>5 </input>
<output>
<ID>OUT</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>8</ID>
<type>AE_OR3</type>
<position>8,-26</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>16 </input>
<input>
<ID>IN_2</ID>15 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>9</ID>
<type>AE_OR3</type>
<position>8,-34</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>13 </input>
<input>
<ID>IN_2</ID>14 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>10</ID>
<type>BA_NAND3</type>
<position>48.5,-8</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>24 </input>
<input>
<ID>IN_2</ID>25 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_AND3</type>
<position>19,-34</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>11 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_REGISTER4</type>
<position>16.5,11.5</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>49 </input>
<input>
<ID>IN_2</ID>48 </input>
<input>
<ID>IN_3</ID>50 </input>
<output>
<ID>OUT_0</ID>61 </output>
<output>
<ID>OUT_1</ID>59 </output>
<output>
<ID>OUT_2</ID>57 </output>
<output>
<ID>OUT_3</ID>55 </output>
<input>
<ID>clear</ID>52 </input>
<input>
<ID>clock</ID>53 </input>
<input>
<ID>count_enable</ID>46 </input>
<input>
<ID>count_up</ID>43 </input>
<input>
<ID>load</ID>45 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>13</ID>
<type>BA_NAND2</type>
<position>48.5,-14</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>BA_NAND2</type>
<position>48.5,-19</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>DE_TO</type>
<position>28.5,-14</position>
<input>
<ID>IN_0</ID>62 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND-OR</lparam></gate>
<gate>
<ID>16</ID>
<type>DE_TO</type>
<position>26,-34</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OR-AND</lparam></gate>
<gate>
<ID>17</ID>
<type>BE_NOR3</type>
<position>48.5,-27</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>35 </input>
<input>
<ID>IN_2</ID>36 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>18</ID>
<type>DA_FROM</type>
<position>2,-6</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A'</lparam></gate>
<gate>
<ID>19</ID>
<type>DA_FROM</type>
<position>2,-8</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B'</lparam></gate>
<gate>
<ID>20</ID>
<type>DA_FROM</type>
<position>2,-10</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C'</lparam></gate>
<gate>
<ID>21</ID>
<type>DA_FROM</type>
<position>2,-13</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C'</lparam></gate>
<gate>
<ID>22</ID>
<type>DA_FROM</type>
<position>2,-15</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D'</lparam></gate>
<gate>
<ID>23</ID>
<type>DA_FROM</type>
<position>2,-18</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>24</ID>
<type>DA_FROM</type>
<position>2,-20</position>
<input>
<ID>IN_0</ID>21 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>25</ID>
<type>DA_FROM</type>
<position>1.5,-24</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>26</ID>
<type>DA_FROM</type>
<position>1.5,-26</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B'</lparam></gate>
<gate>
<ID>27</ID>
<type>DA_FROM</type>
<position>1.5,-28</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D'</lparam></gate>
<gate>
<ID>28</ID>
<type>DA_FROM</type>
<position>1.5,-32</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A'</lparam></gate>
<gate>
<ID>29</ID>
<type>DA_FROM</type>
<position>1.5,-34</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>30</ID>
<type>DA_FROM</type>
<position>1.5,-36</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D'</lparam></gate>
<gate>
<ID>31</ID>
<type>DA_FROM</type>
<position>10,-40</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C'</lparam></gate>
<gate>
<ID>32</ID>
<type>BE_NOR3</type>
<position>48.5,-35</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>38 </input>
<input>
<ID>IN_2</ID>39 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>36</ID>
<type>DD_KEYPAD_HEX</type>
<position>5,12</position>
<output>
<ID>OUT_0</ID>51 </output>
<output>
<ID>OUT_1</ID>49 </output>
<output>
<ID>OUT_2</ID>48 </output>
<output>
<ID>OUT_3</ID>50 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 6</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_TOGGLE</type>
<position>11,18</position>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>39</ID>
<type>DE_TO</type>
<position>68.5,-14</position>
<input>
<ID>IN_0</ID>22 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NAND-NANDX</lparam></gate>
<gate>
<ID>40</ID>
<type>DA_FROM</type>
<position>42,-6</position>
<input>
<ID>IN_0</ID>23 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A'</lparam></gate>
<gate>
<ID>41</ID>
<type>DA_FROM</type>
<position>42,-8</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B'</lparam></gate>
<gate>
<ID>42</ID>
<type>DA_FROM</type>
<position>42,-10</position>
<input>
<ID>IN_0</ID>25 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C'</lparam></gate>
<gate>
<ID>43</ID>
<type>DA_FROM</type>
<position>42,-13</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C'</lparam></gate>
<gate>
<ID>44</ID>
<type>DA_FROM</type>
<position>42,-15</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D'</lparam></gate>
<gate>
<ID>45</ID>
<type>DA_FROM</type>
<position>42,-18</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>46</ID>
<type>DA_FROM</type>
<position>42,-20</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_TOGGLE</type>
<position>17.5,24</position>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>51</ID>
<type>DE_TO</type>
<position>66.5,-35</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NOR-NORX</lparam></gate>
<gate>
<ID>52</ID>
<type>DA_FROM</type>
<position>42,-25</position>
<input>
<ID>IN_0</ID>34 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>53</ID>
<type>DA_FROM</type>
<position>42,-27</position>
<input>
<ID>IN_0</ID>35 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B'</lparam></gate>
<gate>
<ID>54</ID>
<type>DA_FROM</type>
<position>42,-29</position>
<input>
<ID>IN_0</ID>36 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D'</lparam></gate>
<gate>
<ID>55</ID>
<type>DA_FROM</type>
<position>42,-33</position>
<input>
<ID>IN_0</ID>37 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A'</lparam></gate>
<gate>
<ID>56</ID>
<type>DA_FROM</type>
<position>42,-35</position>
<input>
<ID>IN_0</ID>38 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>57</ID>
<type>DA_FROM</type>
<position>42,-37</position>
<input>
<ID>IN_0</ID>39 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D'</lparam></gate>
<gate>
<ID>58</ID>
<type>DA_FROM</type>
<position>50.5,-41</position>
<input>
<ID>IN_0</ID>42 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_TOGGLE</type>
<position>11,21</position>
<output>
<ID>OUT_0</ID>46 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_TOGGLE</type>
<position>23,-2</position>
<output>
<ID>OUT_0</ID>52 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>64</ID>
<type>BB_CLOCK</type>
<position>6.5,2.5</position>
<output>
<ID>CLK</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>66</ID>
<type>DE_TO</type>
<position>31.5,21</position>
<input>
<ID>IN_0</ID>55 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>68</ID>
<type>AE_SMALL_INVERTER</type>
<position>26.5,18</position>
<input>
<ID>IN_0</ID>55 </input>
<output>
<ID>OUT_0</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>69</ID>
<type>DE_TO</type>
<position>31.5,18</position>
<input>
<ID>IN_0</ID>54 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A'</lparam></gate>
<gate>
<ID>70</ID>
<type>DE_TO</type>
<position>31.5,15.5</position>
<input>
<ID>IN_0</ID>57 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>71</ID>
<type>AE_SMALL_INVERTER</type>
<position>26.5,12.5</position>
<input>
<ID>IN_0</ID>57 </input>
<output>
<ID>OUT_0</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>72</ID>
<type>DE_TO</type>
<position>31.5,12.5</position>
<input>
<ID>IN_0</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B'</lparam></gate>
<gate>
<ID>73</ID>
<type>DE_TO</type>
<position>31.5,10</position>
<input>
<ID>IN_0</ID>59 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>74</ID>
<type>AE_SMALL_INVERTER</type>
<position>26.5,7</position>
<input>
<ID>IN_0</ID>59 </input>
<output>
<ID>OUT_0</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>75</ID>
<type>DE_TO</type>
<position>31.5,7</position>
<input>
<ID>IN_0</ID>58 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C'</lparam></gate>
<gate>
<ID>76</ID>
<type>DE_TO</type>
<position>31.5,4</position>
<input>
<ID>IN_0</ID>61 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>77</ID>
<type>AE_SMALL_INVERTER</type>
<position>26.5,1</position>
<input>
<ID>IN_0</ID>61 </input>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>78</ID>
<type>DE_TO</type>
<position>31.5,1</position>
<input>
<ID>IN_0</ID>60 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D'</lparam></gate>
<gate>
<ID>80</ID>
<type>GA_LED</type>
<position>26.5,-10.5</position>
<input>
<ID>N_in2</ID>62 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>GA_LED</type>
<position>24,-31</position>
<input>
<ID>N_in2</ID>2 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>GA_LED</type>
<position>66.5,-11</position>
<input>
<ID>N_in2</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>83</ID>
<type>GA_LED</type>
<position>64.5,-32</position>
<input>
<ID>N_in2</ID>33 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-34,24,-34</points>
<connection>
<GID>11</GID>
<name>OUT</name></connection>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>24 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>24,-34,24,-32</points>
<connection>
<GID>81</GID>
<name>N_in2</name></connection>
<intersection>-34 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-12,15,-8</points>
<intersection>-12 1</intersection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-12,19,-12</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>15 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-8,15,-8</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11.5,-14,19,-14</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<connection>
<GID>7</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-16,19,-16</points>
<connection>
<GID>7</GID>
<name>IN_2</name></connection>
<intersection>15 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>15,-19,15,-16</points>
<intersection>-19 5</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>11,-19,15,-19</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<intersection>15 4</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,-32,13.5,-26</points>
<intersection>-32 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13.5,-32,16,-32</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>13.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-26,13.5,-26</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<intersection>13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11,-34,16,-34</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<connection>
<GID>11</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-6,5.5,-6</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>18</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-13,5.5,-13</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<connection>
<GID>21</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-24,5,-24</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<connection>
<GID>25</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,-40,13.5,-36</points>
<intersection>-40 2</intersection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13.5,-36,16,-36</points>
<connection>
<GID>11</GID>
<name>IN_2</name></connection>
<intersection>13.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12,-40,13.5,-40</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-32,5,-32</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<connection>
<GID>28</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-34,5,-34</points>
<connection>
<GID>9</GID>
<name>IN_1</name></connection>
<connection>
<GID>29</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-36,5,-36</points>
<connection>
<GID>9</GID>
<name>IN_2</name></connection>
<connection>
<GID>30</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-28,5,-28</points>
<connection>
<GID>8</GID>
<name>IN_2</name></connection>
<connection>
<GID>27</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-26,5,-26</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<connection>
<GID>26</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-8,5.5,-8</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<connection>
<GID>19</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-10,5.5,-10</points>
<connection>
<GID>2</GID>
<name>IN_2</name></connection>
<connection>
<GID>20</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-15,5.5,-15</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<connection>
<GID>22</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-18,5,-18</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<connection>
<GID>23</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,-20,5,-20</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<connection>
<GID>24</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>65,-14,66.5,-14</points>
<connection>
<GID>3</GID>
<name>OUT</name></connection>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>66.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>66.5,-14,66.5,-12</points>
<connection>
<GID>82</GID>
<name>N_in2</name></connection>
<intersection>-14 1</intersection></vsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-6,45.5,-6</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<connection>
<GID>10</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-8,45.5,-8</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<connection>
<GID>10</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-10,45.5,-10</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<connection>
<GID>10</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-13,45.5,-13</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<connection>
<GID>13</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-15,45.5,-15</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<connection>
<GID>13</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-18,45.5,-18</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<connection>
<GID>14</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-20,45.5,-20</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<connection>
<GID>14</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-19,55,-16</points>
<intersection>-19 2</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-16,59,-16</points>
<connection>
<GID>3</GID>
<name>IN_2</name></connection>
<intersection>55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-19,55,-19</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51.5,-14,59,-14</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<connection>
<GID>13</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-12,55,-8</points>
<intersection>-12 1</intersection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-12,59,-12</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-8,55,-8</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>63,-35,64.5,-35</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>64.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>64.5,-35,64.5,-33</points>
<connection>
<GID>83</GID>
<name>N_in2</name></connection>
<intersection>-35 1</intersection></vsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-25,45.5,-25</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<connection>
<GID>17</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-27,45.5,-27</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<connection>
<GID>17</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-29,45.5,-29</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<connection>
<GID>17</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-33,45.5,-33</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<connection>
<GID>32</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-35,45.5,-35</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<connection>
<GID>32</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-37,45.5,-37</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<connection>
<GID>32</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-33,54,-27</points>
<intersection>-33 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-33,57,-33</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-27,54,-27</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51.5,-35,57,-35</points>
<connection>
<GID>32</GID>
<name>OUT</name></connection>
<connection>
<GID>6</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-41,54.5,-37</points>
<intersection>-41 2</intersection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-37,57,-37</points>
<connection>
<GID>6</GID>
<name>IN_2</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52.5,-41,54.5,-41</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,16.5,17.5,22</points>
<connection>
<GID>12</GID>
<name>count_up</name></connection>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,16.5,15.5,18</points>
<connection>
<GID>12</GID>
<name>load</name></connection>
<intersection>18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,18,15.5,18</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,16.5,16.5,21</points>
<connection>
<GID>12</GID>
<name>count_enable</name></connection>
<intersection>21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,21,16.5,21</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<intersection>16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,12.5,11.5,13</points>
<intersection>12.5 1</intersection>
<intersection>13 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11.5,12.5,12.5,12.5</points>
<connection>
<GID>12</GID>
<name>IN_2</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10,13,11.5,13</points>
<connection>
<GID>36</GID>
<name>OUT_2</name></connection>
<intersection>11.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,11,11.5,11.5</points>
<intersection>11 2</intersection>
<intersection>11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11.5,11.5,12.5,11.5</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10,11,11.5,11</points>
<connection>
<GID>36</GID>
<name>OUT_1</name></connection>
<intersection>11.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,13.5,11.5,15</points>
<intersection>13.5 1</intersection>
<intersection>15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11.5,13.5,12.5,13.5</points>
<connection>
<GID>12</GID>
<name>IN_3</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10,15,11.5,15</points>
<connection>
<GID>36</GID>
<name>OUT_3</name></connection>
<intersection>11.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,9,11.5,10.5</points>
<intersection>9 2</intersection>
<intersection>10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11.5,10.5,12.5,10.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10,9,11.5,9</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>11.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-2,17.5,7.5</points>
<connection>
<GID>12</GID>
<name>clear</name></connection>
<intersection>-2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-2,21,-2</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,2.5,15.5,7.5</points>
<connection>
<GID>12</GID>
<name>clock</name></connection>
<intersection>2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10.5,2.5,15.5,2.5</points>
<connection>
<GID>64</GID>
<name>CLK</name></connection>
<intersection>15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,18,29.5,18</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,13.5,23,21</points>
<intersection>13.5 6</intersection>
<intersection>18 2</intersection>
<intersection>21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,21,29.5,21</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,18,24.5,18</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>20.5,13.5,23,13.5</points>
<connection>
<GID>12</GID>
<name>OUT_3</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,12.5,29.5,12.5</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,12.5,24.5,15.5</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>12.5 4</intersection>
<intersection>15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,15.5,29.5,15.5</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>20.5,12.5,24.5,12.5</points>
<connection>
<GID>12</GID>
<name>OUT_2</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>13</ID>
<points>28.5,7,29.5,7</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,7,24.5,11.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>10 1</intersection>
<intersection>11.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,10,29.5,10</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>20.5,11.5,24.5,11.5</points>
<connection>
<GID>12</GID>
<name>OUT_1</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,1,29.5,1</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,1,23,10.5</points>
<intersection>1 2</intersection>
<intersection>4 1</intersection>
<intersection>10.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,4,29.5,4</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,1,24.5,1</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>20.5,10.5,23,10.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-14,26.5,-11.5</points>
<connection>
<GID>80</GID>
<name>N_in2</name></connection>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-14,26.5,-14</points>
<connection>
<GID>7</GID>
<name>OUT</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,116.147,1079.94,-502.863</PageViewport></page 1>
<page 2>
<PageViewport>0,116.147,1079.94,-502.863</PageViewport></page 2>
<page 3>
<PageViewport>0,116.147,1079.94,-502.863</PageViewport></page 3>
<page 4>
<PageViewport>0,116.147,1079.94,-502.863</PageViewport></page 4>
<page 5>
<PageViewport>0,116.147,1079.94,-502.863</PageViewport></page 5>
<page 6>
<PageViewport>0,116.147,1079.94,-502.863</PageViewport></page 6>
<page 7>
<PageViewport>0,116.147,1079.94,-502.863</PageViewport></page 7>
<page 8>
<PageViewport>0,116.147,1079.94,-502.863</PageViewport></page 8>
<page 9>
<PageViewport>0,116.147,1079.94,-502.863</PageViewport></page 9></circuit>