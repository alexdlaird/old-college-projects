<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-40.275,6.93531,59.775,-50.4123</PageViewport>
<gate>
<ID>1</ID>
<type>AE_REGISTER8</type>
<position>29.5,-26.5</position>
<output>
<ID>OUT_0</ID>53 </output>
<output>
<ID>OUT_1</ID>54 </output>
<output>
<ID>OUT_2</ID>55 </output>
<output>
<ID>OUT_3</ID>56 </output>
<input>
<ID>clear</ID>59 </input>
<input>
<ID>clock</ID>48 </input>
<input>
<ID>count_enable</ID>6 </input>
<input>
<ID>count_up</ID>6 </input>
<input>
<ID>load</ID>10 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 10</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>15,-7.5</position>
<gparam>LABEL_TEXT X(input)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>DD_KEYPAD_HEX</type>
<position>-21.5,-7.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<output>
<ID>OUT_1</ID>2 </output>
<output>
<ID>OUT_2</ID>3 </output>
<output>
<ID>OUT_3</ID>4 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 2</lparam></gate>
<gate>
<ID>4</ID>
<type>FF_GND</type>
<position>-23.5,-21</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>5</ID>
<type>DA_FROM</type>
<position>-19.5,-31</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Not_Done</lparam></gate>
<gate>
<ID>6</ID>
<type>AE_SMALL_INVERTER</type>
<position>35,-22.5</position>
<input>
<ID>IN_0</ID>57 </input>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7</ID>
<type>GF_LED_DISPLAY_4BIT_OUT</type>
<position>-11.5,-8</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>3 </input>
<input>
<ID>IN_3</ID>4 </input>
<output>
<ID>OUT_0</ID>17 </output>
<output>
<ID>OUT_1</ID>15 </output>
<output>
<ID>OUT_2</ID>14 </output>
<output>
<ID>OUT_3</ID>16 </output>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>8</ID>
<type>DD_KEYPAD_HEX</type>
<position>0,-7.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<output>
<ID>OUT_1</ID>8 </output>
<output>
<ID>OUT_2</ID>19 </output>
<output>
<ID>OUT_3</ID>21 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 10</lparam></gate>
<gate>
<ID>9</ID>
<type>GF_LED_DISPLAY_4BIT_OUT</type>
<position>10,-8</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>8 </input>
<input>
<ID>IN_2</ID>19 </input>
<input>
<ID>IN_3</ID>21 </input>
<output>
<ID>OUT_0</ID>49 </output>
<output>
<ID>OUT_1</ID>50 </output>
<output>
<ID>OUT_2</ID>51 </output>
<output>
<ID>OUT_3</ID>52 </output>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 10</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>10</ID>
<type>FF_GND</type>
<position>25,-20.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>11</ID>
<type>GA_LED</type>
<position>27,-3</position>
<input>
<ID>N_in0</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>DE_TO</type>
<position>39,-19.5</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Not_Done</lparam></gate>
<gate>
<ID>13</ID>
<type>DE_TO</type>
<position>39,-24.5</position>
<input>
<ID>IN_0</ID>57 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Done</lparam></gate>
<gate>
<ID>14</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-15,-25.5</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>43 </input>
<input>
<ID>IN_2</ID>42 </input>
<input>
<ID>IN_3</ID>41 </input>
<input>
<ID>IN_B_0</ID>17 </input>
<input>
<ID>IN_B_1</ID>15 </input>
<input>
<ID>IN_B_2</ID>14 </input>
<input>
<ID>IN_B_3</ID>16 </input>
<output>
<ID>OUT_0</ID>33 </output>
<output>
<ID>OUT_1</ID>32 </output>
<output>
<ID>OUT_2</ID>31 </output>
<output>
<ID>OUT_3</ID>30 </output>
<input>
<ID>carry_in</ID>18 </input>
<output>
<ID>carry_out</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_TOGGLE</type>
<position>9.5,1.5</position>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>30.5,-7</position>
<gparam>LABEL_TEXT Alex Laird</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>DA_FROM</type>
<position>25,-33</position>
<input>
<ID>IN_0</ID>48 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>18</ID>
<type>DA_FROM</type>
<position>23,-3</position>
<input>
<ID>IN_0</ID>23 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Done</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>-31,-18.5</position>
<gparam>LABEL_TEXT 8bit Full Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>DE_TO</type>
<position>-26,-44</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>22</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>47.5,-34.5</position>
<output>
<ID>A_equal_B</ID>57 </output>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>54 </input>
<input>
<ID>IN_2</ID>55 </input>
<input>
<ID>IN_3</ID>56 </input>
<input>
<ID>IN_B_0</ID>49 </input>
<input>
<ID>IN_B_1</ID>50 </input>
<input>
<ID>IN_B_2</ID>51 </input>
<input>
<ID>IN_B_3</ID>52 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>-25.5,-38.5</position>
<gparam>LABEL_TEXT Accumulator</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-32,-25.5</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>12 </input>
<input>
<ID>IN_2</ID>20 </input>
<input>
<ID>IN_3</ID>22 </input>
<input>
<ID>IN_B_0</ID>9 </input>
<input>
<ID>IN_B_1</ID>9 </input>
<input>
<ID>IN_B_2</ID>9 </input>
<input>
<ID>IN_B_3</ID>9 </input>
<output>
<ID>OUT_0</ID>29 </output>
<output>
<ID>OUT_1</ID>28 </output>
<output>
<ID>OUT_2</ID>27 </output>
<output>
<ID>OUT_3</ID>26 </output>
<input>
<ID>carry_in</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>26</ID>
<type>FF_GND</type>
<position>-4.5,-25.5</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>30</ID>
<type>DA_FROM</type>
<position>27,-36</position>
<input>
<ID>IN_0</ID>59 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Load/Mult</lparam></gate>
<gate>
<ID>35</ID>
<type>DE_TO</type>
<position>15,1.5</position>
<input>
<ID>IN_0</ID>36 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Load/Mult</lparam></gate>
<gate>
<ID>38</ID>
<type>AE_REGISTER8</type>
<position>-6,-37</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>32 </input>
<input>
<ID>IN_2</ID>31 </input>
<input>
<ID>IN_3</ID>30 </input>
<input>
<ID>IN_4</ID>29 </input>
<input>
<ID>IN_5</ID>28 </input>
<input>
<ID>IN_6</ID>27 </input>
<input>
<ID>IN_7</ID>26 </input>
<output>
<ID>OUT_0</ID>44 </output>
<output>
<ID>OUT_1</ID>43 </output>
<output>
<ID>OUT_2</ID>42 </output>
<output>
<ID>OUT_3</ID>41 </output>
<output>
<ID>OUT_4</ID>11 </output>
<output>
<ID>OUT_5</ID>12 </output>
<output>
<ID>OUT_6</ID>20 </output>
<output>
<ID>OUT_7</ID>22 </output>
<output>
<ID>carry_out</ID>39 </output>
<input>
<ID>clear</ID>35 </input>
<input>
<ID>clock</ID>34 </input>
<input>
<ID>count_enable</ID>40 </input>
<input>
<ID>count_up</ID>40 </input>
<input>
<ID>load</ID>5 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 20</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>42</ID>
<type>DA_FROM</type>
<position>-9,-43.5</position>
<input>
<ID>IN_0</ID>34 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>44</ID>
<type>DA_FROM</type>
<position>-9,-45.5</position>
<input>
<ID>IN_0</ID>35 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Load/Mult</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>-38.5,2</position>
<gparam>LABEL_TEXT 4bit Repeated Addition Mulitplier</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>GA_LED</type>
<position>-0.5,-30.5</position>
<input>
<ID>N_in0</ID>39 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>BB_CLOCK</type>
<position>-33,-44</position>
<output>
<ID>CLK</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>50</ID>
<type>FF_GND</type>
<position>1.5,-29.5</position>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>52</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>12,-37</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>43 </input>
<input>
<ID>IN_2</ID>42 </input>
<input>
<ID>IN_3</ID>41 </input>
<input>
<ID>IN_4</ID>11 </input>
<input>
<ID>IN_5</ID>12 </input>
<input>
<ID>IN_6</ID>20 </input>
<input>
<ID>IN_7</ID>22 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 20</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15.5,-10.5,-15.5,-9</points>
<intersection>-10.5 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15.5,-9,-14.5,-9</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-16.5,-10.5,-15.5,-10.5</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>-15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15.5,-8.5,-15.5,-8</points>
<intersection>-8.5 2</intersection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15.5,-8,-14.5,-8</points>
<connection>
<GID>7</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-16.5,-8.5,-15.5,-8.5</points>
<connection>
<GID>3</GID>
<name>OUT_1</name></connection>
<intersection>-15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15.5,-7,-15.5,-6.5</points>
<intersection>-7 2</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16.5,-6.5,-15.5,-6.5</points>
<connection>
<GID>3</GID>
<name>OUT_2</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-15.5,-7,-14.5,-7</points>
<connection>
<GID>7</GID>
<name>IN_2</name></connection>
<intersection>-15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15.5,-6,-15.5,-4.5</points>
<intersection>-6 2</intersection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16.5,-4.5,-15.5,-4.5</points>
<connection>
<GID>3</GID>
<name>OUT_3</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-15.5,-6,-14.5,-6</points>
<connection>
<GID>7</GID>
<name>IN_3</name></connection>
<intersection>-15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-17.5,-31,-7,-31</points>
<connection>
<GID>38</GID>
<name>load</name></connection>
<connection>
<GID>5</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>29.5,-19.5,37,-19.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>29.5 12</intersection>
<intersection>30.5 13</intersection>
<intersection>35 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>35,-20.5,35,-19.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>-19.5 3</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>29.5,-20.5,29.5,-19.5</points>
<connection>
<GID>1</GID>
<name>count_enable</name></connection>
<intersection>-19.5 3</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>30.5,-20.5,30.5,-19.5</points>
<connection>
<GID>1</GID>
<name>count_up</name></connection>
<intersection>-19.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-10.5,6,-9</points>
<intersection>-10.5 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6,-9,7,-9</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5,-10.5,6,-10.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-8.5,6,-8</points>
<intersection>-8.5 2</intersection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6,-8,7,-8</points>
<connection>
<GID>9</GID>
<name>IN_1</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5,-8.5,6,-8.5</points>
<connection>
<GID>8</GID>
<name>OUT_1</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-27,-21.5,-27,-20</points>
<connection>
<GID>24</GID>
<name>IN_B_0</name></connection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-30,-20,-23.5,-20</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-30 6</intersection>
<intersection>-29 7</intersection>
<intersection>-28 8</intersection>
<intersection>-27 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-30,-21.5,-30,-20</points>
<connection>
<GID>24</GID>
<name>IN_B_3</name></connection>
<intersection>-20 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-29,-21.5,-29,-20</points>
<connection>
<GID>24</GID>
<name>IN_B_2</name></connection>
<intersection>-20 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-28,-21.5,-28,-20</points>
<connection>
<GID>24</GID>
<name>IN_B_1</name></connection>
<intersection>-20 2</intersection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>25,-18.5,28.5,-18.5</points>
<intersection>25 3</intersection>
<intersection>28.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25,-19.5,25,-18.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>-18.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>28.5,-20.5,28.5,-18.5</points>
<connection>
<GID>1</GID>
<name>load</name></connection>
<intersection>-18.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-21.5,-34,-16</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34,-16,5,-16</points>
<intersection>-34 0</intersection>
<intersection>5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>5,-36,5,-16</points>
<intersection>-36 3</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-2,-36,7,-36</points>
<connection>
<GID>38</GID>
<name>OUT_4</name></connection>
<connection>
<GID>52</GID>
<name>IN_4</name></connection>
<intersection>5 2</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-35,-15.5,5.5,-15.5</points>
<intersection>-35 3</intersection>
<intersection>5.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-35,-21.5,-35,-15.5</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>-15.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>5.5,-35,5.5,-15.5</points>
<intersection>-35 6</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-2,-35,7,-35</points>
<connection>
<GID>38</GID>
<name>OUT_5</name></connection>
<connection>
<GID>52</GID>
<name>IN_5</name></connection>
<intersection>5.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-24,-24.5,-23,-24.5</points>
<connection>
<GID>14</GID>
<name>carry_out</name></connection>
<connection>
<GID>24</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-21.5,-12,-12</points>
<connection>
<GID>14</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>7</GID>
<name>OUT_2</name></connection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,-21.5,-11,-12</points>
<connection>
<GID>14</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>7</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13,-21.5,-13,-12</points>
<connection>
<GID>14</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>7</GID>
<name>OUT_3</name></connection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,-21.5,-10,-12</points>
<connection>
<GID>14</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-7,-24.5,-4.5,-24.5</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<connection>
<GID>14</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-7,6,-6.5</points>
<intersection>-7 2</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,-6.5,6,-6.5</points>
<connection>
<GID>8</GID>
<name>OUT_2</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6,-7,7,-7</points>
<connection>
<GID>9</GID>
<name>IN_2</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-36,-15,6,-15</points>
<intersection>-36 3</intersection>
<intersection>6 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-36,-21.5,-36,-15</points>
<connection>
<GID>24</GID>
<name>IN_2</name></connection>
<intersection>-15 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>6,-34,6,-15</points>
<intersection>-34 6</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-2,-34,7,-34</points>
<connection>
<GID>38</GID>
<name>OUT_6</name></connection>
<connection>
<GID>52</GID>
<name>IN_6</name></connection>
<intersection>6 4</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-6,6,-4.5</points>
<intersection>-6 2</intersection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,-4.5,6,-4.5</points>
<connection>
<GID>8</GID>
<name>OUT_3</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6,-6,7,-6</points>
<connection>
<GID>9</GID>
<name>IN_3</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-37,-14.5,6.5,-14.5</points>
<intersection>-37 3</intersection>
<intersection>6.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-37,-21.5,-37,-14.5</points>
<connection>
<GID>24</GID>
<name>IN_3</name></connection>
<intersection>-14.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>6.5,-33,6.5,-14.5</points>
<intersection>-33 6</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-2,-33,7,-33</points>
<connection>
<GID>38</GID>
<name>OUT_7</name></connection>
<connection>
<GID>52</GID>
<name>IN_7</name></connection>
<intersection>6.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25,-3,26,-3</points>
<connection>
<GID>11</GID>
<name>N_in0</name></connection>
<connection>
<GID>18</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-29,-44,-28,-44</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<connection>
<GID>49</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33.5,-33,-33.5,-29.5</points>
<connection>
<GID>24</GID>
<name>OUT_3</name></connection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-33.5,-33,-10,-33</points>
<connection>
<GID>38</GID>
<name>IN_7</name></connection>
<intersection>-33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32.5,-34,-32.5,-29.5</points>
<connection>
<GID>24</GID>
<name>OUT_2</name></connection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-32.5,-34,-10,-34</points>
<connection>
<GID>38</GID>
<name>IN_6</name></connection>
<intersection>-32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-31.5,-35,-31.5,-29.5</points>
<connection>
<GID>24</GID>
<name>OUT_1</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-31.5,-35,-10,-35</points>
<connection>
<GID>38</GID>
<name>IN_5</name></connection>
<intersection>-31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30.5,-36,-30.5,-29.5</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-30.5,-36,-10,-36</points>
<connection>
<GID>38</GID>
<name>IN_4</name></connection>
<intersection>-30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-37,-16.5,-29.5</points>
<connection>
<GID>14</GID>
<name>OUT_3</name></connection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16.5,-37,-10,-37</points>
<connection>
<GID>38</GID>
<name>IN_3</name></connection>
<intersection>-16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15.5,-38,-15.5,-29.5</points>
<connection>
<GID>14</GID>
<name>OUT_2</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15.5,-38,-10,-38</points>
<connection>
<GID>38</GID>
<name>IN_2</name></connection>
<intersection>-15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-39,-14.5,-29.5</points>
<connection>
<GID>14</GID>
<name>OUT_1</name></connection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,-39,-10,-39</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,-40,-13.5,-29.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13.5,-40,-10,-40</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>-13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7,-43.5,-7,-42</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<connection>
<GID>38</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-45.5,-5,-42</points>
<connection>
<GID>38</GID>
<name>clear</name></connection>
<intersection>-45.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7,-45.5,-5,-45.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>-5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11.5,1.5,13,1.5</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<intersection>13 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>13,1.5,13,1.5</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>1.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-31,-4,-30.5</points>
<connection>
<GID>38</GID>
<name>carry_out</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4,-30.5,-1.5,-30.5</points>
<connection>
<GID>48</GID>
<name>N_in0</name></connection>
<intersection>-4 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-31,-5,-28.5</points>
<connection>
<GID>38</GID>
<name>count_up</name></connection>
<intersection>-31 4</intersection>
<intersection>-28.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-5,-28.5,1.5,-28.5</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>-5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-6,-31,-5,-31</points>
<connection>
<GID>38</GID>
<name>count_enable</name></connection>
<intersection>-5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-37,7,-37</points>
<connection>
<GID>38</GID>
<name>OUT_3</name></connection>
<connection>
<GID>52</GID>
<name>IN_3</name></connection>
<intersection>4 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>4,-37,4,-17</points>
<intersection>-37 1</intersection>
<intersection>-17 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-20,-17,4,-17</points>
<intersection>-20 9</intersection>
<intersection>4 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-20,-21.5,-20,-17</points>
<connection>
<GID>14</GID>
<name>IN_3</name></connection>
<intersection>-17 8</intersection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-38,7,-38</points>
<connection>
<GID>38</GID>
<name>OUT_2</name></connection>
<connection>
<GID>52</GID>
<name>IN_2</name></connection>
<intersection>3.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>3.5,-38,3.5,-17.5</points>
<intersection>-38 1</intersection>
<intersection>-17.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-19,-17.5,3.5,-17.5</points>
<intersection>-19 9</intersection>
<intersection>3.5 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-19,-21.5,-19,-17.5</points>
<connection>
<GID>14</GID>
<name>IN_2</name></connection>
<intersection>-17.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-39,7,-39</points>
<connection>
<GID>38</GID>
<name>OUT_1</name></connection>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>3 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>3,-39,3,-18</points>
<intersection>-39 1</intersection>
<intersection>-18 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-18,-18,3,-18</points>
<intersection>-18 9</intersection>
<intersection>3 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-18,-21.5,-18,-18</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>-18 8</intersection></vsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-40,7,-40</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>2.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>2.5,-40,2.5,-18.5</points>
<intersection>-40 1</intersection>
<intersection>-18.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-17,-18.5,2.5,-18.5</points>
<intersection>-17 9</intersection>
<intersection>2.5 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-17,-21.5,-17,-18.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>-18.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-33,28.5,-31.5</points>
<connection>
<GID>1</GID>
<name>clock</name></connection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-33,28.5,-33</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-30.5,52.5,-15</points>
<connection>
<GID>22</GID>
<name>IN_B_0</name></connection>
<intersection>-15 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>11.5,-15,11.5,-12</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-15,52.5,-15</points>
<intersection>11.5 1</intersection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-30.5,51.5,-15.5</points>
<connection>
<GID>22</GID>
<name>IN_B_1</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>10.5,-15.5,10.5,-12</points>
<connection>
<GID>9</GID>
<name>OUT_1</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>10.5,-15.5,51.5,-15.5</points>
<intersection>10.5 1</intersection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-30.5,50.5,-16</points>
<connection>
<GID>22</GID>
<name>IN_B_2</name></connection>
<intersection>-16 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>9.5,-16,9.5,-12</points>
<connection>
<GID>9</GID>
<name>OUT_2</name></connection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>9.5,-16,50.5,-16</points>
<intersection>9.5 1</intersection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-30.5,49.5,-16.5</points>
<connection>
<GID>22</GID>
<name>IN_B_3</name></connection>
<intersection>-16.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>8.5,-16.5,8.5,-12</points>
<connection>
<GID>9</GID>
<name>OUT_3</name></connection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-16.5,49.5,-16.5</points>
<intersection>8.5 1</intersection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-30.5,45.5,-29.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-29.5,45.5,-29.5</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-30.5,44.5,-28.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-28.5,44.5,-28.5</points>
<connection>
<GID>1</GID>
<name>OUT_1</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-30.5,43.5,-27.5</points>
<connection>
<GID>22</GID>
<name>IN_2</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-27.5,43.5,-27.5</points>
<connection>
<GID>1</GID>
<name>OUT_2</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-30.5,42.5,-26.5</points>
<connection>
<GID>22</GID>
<name>IN_3</name></connection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-26.5,42.5,-26.5</points>
<connection>
<GID>1</GID>
<name>OUT_3</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-34.5,35,-24.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>-34.5 1</intersection>
<intersection>-24.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-34.5,39.5,-34.5</points>
<connection>
<GID>22</GID>
<name>A_equal_B</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-24.5,37,-24.5</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-36,30.5,-31.5</points>
<connection>
<GID>1</GID>
<name>clear</name></connection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-36,30.5,-36</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>99.7449,-15.1565,150.791,-44.4156</PageViewport></page 1>
<page 2>
<PageViewport>-4.36369,198.478,1293.64,-545.522</PageViewport></page 2>
<page 3>
<PageViewport>-4.36369,198.478,1293.64,-545.522</PageViewport></page 3>
<page 4>
<PageViewport>-4.36369,198.478,1293.64,-545.522</PageViewport></page 4>
<page 5>
<PageViewport>-4.36369,198.478,1293.64,-545.522</PageViewport></page 5>
<page 6>
<PageViewport>-4.36369,198.478,1293.64,-545.522</PageViewport></page 6>
<page 7>
<PageViewport>-4.36369,198.478,1293.64,-545.522</PageViewport></page 7>
<page 8>
<PageViewport>-4.36369,198.478,1293.64,-545.522</PageViewport></page 8>
<page 9>
<PageViewport>-4.36369,198.478,1293.64,-545.522</PageViewport></page 9></circuit>