<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-44.1375,8.773,25.6875,-31.25</PageViewport>
<gate>
<ID>2</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>18,2.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>2 </input>
<input>
<ID>IN_3</ID>1 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>6</ID>
<type>DA_FROM</type>
<position>11,6</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 0.3</lparam></gate>
<gate>
<ID>7</ID>
<type>DA_FROM</type>
<position>11,4</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 0.2</lparam></gate>
<gate>
<ID>8</ID>
<type>DA_FROM</type>
<position>11,2</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 0.1</lparam></gate>
<gate>
<ID>9</ID>
<type>DA_FROM</type>
<position>11,0</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 0.0</lparam></gate>
<gate>
<ID>10</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>18,-7</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>6 </input>
<input>
<ID>IN_3</ID>5 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>11</ID>
<type>DA_FROM</type>
<position>11,-3.5</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1.3</lparam></gate>
<gate>
<ID>12</ID>
<type>DA_FROM</type>
<position>11,-5.5</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1.2</lparam></gate>
<gate>
<ID>13</ID>
<type>DA_FROM</type>
<position>11,-7.5</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1.1</lparam></gate>
<gate>
<ID>14</ID>
<type>DA_FROM</type>
<position>11,-9.5</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1.0</lparam></gate>
<gate>
<ID>15</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>18,-16.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>11 </input>
<input>
<ID>IN_2</ID>10 </input>
<input>
<ID>IN_3</ID>9 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>16</ID>
<type>DA_FROM</type>
<position>11,-13</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 2.3</lparam></gate>
<gate>
<ID>17</ID>
<type>DA_FROM</type>
<position>11,-15</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 2.2</lparam></gate>
<gate>
<ID>18</ID>
<type>DA_FROM</type>
<position>11,-17</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 2.1</lparam></gate>
<gate>
<ID>19</ID>
<type>DA_FROM</type>
<position>11,-19</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 2.0</lparam></gate>
<gate>
<ID>20</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>18,-26</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>15 </input>
<input>
<ID>IN_2</ID>14 </input>
<input>
<ID>IN_3</ID>13 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>21</ID>
<type>DA_FROM</type>
<position>11,-22.5</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 3.3</lparam></gate>
<gate>
<ID>22</ID>
<type>DA_FROM</type>
<position>11,-24.5</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 3.2</lparam></gate>
<gate>
<ID>23</ID>
<type>DA_FROM</type>
<position>11,-26.5</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 3.1</lparam></gate>
<gate>
<ID>24</ID>
<type>DA_FROM</type>
<position>11,-28.5</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 3.0</lparam></gate>
<gate>
<ID>26</ID>
<type>BE_TRI_STATE_LOW</type>
<position>-22,-4</position>
<input>
<ID>ENABLE_0</ID>29 </input>
<input>
<ID>IN_0</ID>21 </input>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>28</ID>
<type>BA_TRI_STATE</type>
<position>-5,-4</position>
<input>
<ID>ENABLE_0</ID>29 </input>
<input>
<ID>IN_0</ID>1019 </input>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>31</ID>
<type>BE_TRI_STATE_LOW</type>
<position>-22,-9</position>
<input>
<ID>ENABLE_0</ID>29 </input>
<input>
<ID>IN_0</ID>22 </input>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>32</ID>
<type>BA_TRI_STATE</type>
<position>-5,-9</position>
<input>
<ID>ENABLE_0</ID>29 </input>
<input>
<ID>IN_0</ID>1020 </input>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>34</ID>
<type>BE_TRI_STATE_LOW</type>
<position>-22,-14</position>
<input>
<ID>ENABLE_0</ID>29 </input>
<input>
<ID>IN_0</ID>23 </input>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>35</ID>
<type>BA_TRI_STATE</type>
<position>-5,-14</position>
<input>
<ID>ENABLE_0</ID>29 </input>
<input>
<ID>IN_0</ID>1021 </input>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>37</ID>
<type>BE_TRI_STATE_LOW</type>
<position>-22,-19</position>
<input>
<ID>ENABLE_0</ID>29 </input>
<input>
<ID>IN_0</ID>24 </input>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>38</ID>
<type>BA_TRI_STATE</type>
<position>-5,-19</position>
<input>
<ID>ENABLE_0</ID>29 </input>
<input>
<ID>IN_0</ID>1022 </input>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>41</ID>
<type>DD_KEYPAD_HEX</type>
<position>-34.5,-11.5</position>
<output>
<ID>OUT_0</ID>24 </output>
<output>
<ID>OUT_1</ID>23 </output>
<output>
<ID>OUT_2</ID>22 </output>
<output>
<ID>OUT_3</ID>21 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 10</lparam></gate>
<gate>
<ID>43</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>-8,4.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>26 </input>
<input>
<ID>IN_2</ID>27 </input>
<input>
<ID>IN_3</ID>28 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 10</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>44</ID>
<type>DE_TO</type>
<position>-10.5,-24</position>
<input>
<ID>IN_0</ID>25 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>45</ID>
<type>DE_TO</type>
<position>-10.5,-26</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>46</ID>
<type>DE_TO</type>
<position>-10.5,-28</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>47</ID>
<type>DE_TO</type>
<position>-10.5,-30</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_TOGGLE</type>
<position>-29,0.5</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>51</ID>
<type>CC_PULSE</type>
<position>-29,4</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_TOGGLE</type>
<position>-29,7.5</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>55</ID>
<type>DE_TO</type>
<position>-24,7.5</position>
<input>
<ID>IN_0</ID>31 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Reset</lparam></gate>
<gate>
<ID>57</ID>
<type>DE_TO</type>
<position>-24,4</position>
<input>
<ID>IN_0</ID>32 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>59</ID>
<type>DE_TO</type>
<position>-0.5,-24</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r/w</lparam></gate>
<gate>
<ID>61</ID>
<type>DE_TO</type>
<position>0.5,-26</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /r/w</lparam></gate>
<gate>
<ID>63</ID>
<type>AE_SMALL_INVERTER</type>
<position>-4.5,-26</position>
<input>
<ID>IN_0</ID>29 </input>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>-36.5,7.5</position>
<gparam>LABEL_TEXT Reset</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>-36,4</position>
<gparam>LABEL_TEXT Clock</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>-35,0.5</position>
<gparam>LABEL_TEXT R/W</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1297</ID>
<type>DA_FROM</type>
<position>1.5,-4</position>
<input>
<ID>IN_0</ID>1019 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID 0.3</lparam></gate>
<gate>
<ID>1298</ID>
<type>DA_FROM</type>
<position>1.5,-9</position>
<input>
<ID>IN_0</ID>1020 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID 0.2</lparam></gate>
<gate>
<ID>1299</ID>
<type>DA_FROM</type>
<position>1.5,-14</position>
<input>
<ID>IN_0</ID>1021 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID 0.1</lparam></gate>
<gate>
<ID>1300</ID>
<type>DA_FROM</type>
<position>1.5,-19</position>
<input>
<ID>IN_0</ID>1022 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID 0.0</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,6,15,6</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>15 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>15,4.5,15,6</points>
<connection>
<GID>2</GID>
<name>IN_3</name></connection>
<intersection>6 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,4,15,4</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>15 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>15,3.5,15,4</points>
<connection>
<GID>2</GID>
<name>IN_2</name></connection>
<intersection>4 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,2,15,2.5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,2,15,2</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,0,15,1.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,0,15,0</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-3.5,15,-3.5</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>15 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>15,-5,15,-3.5</points>
<connection>
<GID>10</GID>
<name>IN_3</name></connection>
<intersection>-3.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-5.5,15,-5.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>15 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>15,-6,15,-5.5</points>
<connection>
<GID>10</GID>
<name>IN_2</name></connection>
<intersection>-5.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-7.5,15,-7</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,-7.5,15,-7.5</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-9.5,15,-8</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,-9.5,15,-9.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-13,15,-13</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>15 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>15,-14.5,15,-13</points>
<connection>
<GID>15</GID>
<name>IN_3</name></connection>
<intersection>-13 1</intersection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-15,15,-15</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>15 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>15,-15.5,15,-15</points>
<connection>
<GID>15</GID>
<name>IN_2</name></connection>
<intersection>-15 1</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-17,15,-16.5</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,-17,15,-17</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-19,15,-17.5</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,-19,15,-19</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-22.5,15,-22.5</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>15 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>15,-24,15,-22.5</points>
<connection>
<GID>20</GID>
<name>IN_3</name></connection>
<intersection>-22.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-24.5,15,-24.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>15 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>15,-25,15,-24.5</points>
<connection>
<GID>20</GID>
<name>IN_2</name></connection>
<intersection>-24.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-26.5,15,-26</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,-26.5,15,-26.5</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-28.5,15,-27</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,-28.5,15,-28.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26.5,-8.5,-26.5,-4</points>
<intersection>-8.5 2</intersection>
<intersection>-4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-26.5,-4,-25,-4</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>-26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-29.5,-8.5,-26.5,-8.5</points>
<connection>
<GID>41</GID>
<name>OUT_3</name></connection>
<intersection>-26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25.5,-10.5,-25.5,-9</points>
<intersection>-10.5 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25.5,-9,-25,-9</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>-25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-29.5,-10.5,-25.5,-10.5</points>
<connection>
<GID>41</GID>
<name>OUT_2</name></connection>
<intersection>-25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25.5,-14,-25.5,-12.5</points>
<intersection>-14 1</intersection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25.5,-14,-25,-14</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>-25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-29.5,-12.5,-25.5,-12.5</points>
<connection>
<GID>41</GID>
<name>OUT_1</name></connection>
<intersection>-25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26.5,-19,-26.5,-14.5</points>
<intersection>-19 1</intersection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-26.5,-19,-25,-19</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>-26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-29.5,-14.5,-26.5,-14.5</points>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection>
<intersection>-26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12.5,-24,-12.5,3.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>-19 3</intersection>
<intersection>3.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-12.5,3.5,-11,3.5</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>-12.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-19.5,-19,-7.5,-19</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>-12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,-26,-14,4.5</points>
<intersection>-26 2</intersection>
<intersection>-14 3</intersection>
<intersection>4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14,4.5,-11,4.5</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-14,-26,-12.5,-26</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-19.5,-14,-7.5,-14</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15.5,-28,-15.5,5.5</points>
<intersection>-28 2</intersection>
<intersection>-9 3</intersection>
<intersection>5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15.5,5.5,-11,5.5</points>
<connection>
<GID>43</GID>
<name>IN_2</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-15.5,-28,-12.5,-28</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-19.5,-9,-7.5,-9</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>-15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-17,-30,-17,6.5</points>
<intersection>-30 1</intersection>
<intersection>-4 3</intersection>
<intersection>6.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-17,-30,-12.5,-30</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>-17 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-17,6.5,-11,6.5</points>
<connection>
<GID>43</GID>
<name>IN_3</name></connection>
<intersection>-17 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-19.5,-4,-7.5,-4</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>-17 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7,-26,-7,-6.5</points>
<intersection>-26 20</intersection>
<intersection>-24 11</intersection>
<intersection>-21.5 1</intersection>
<intersection>-16.5 22</intersection>
<intersection>-11.5 24</intersection>
<intersection>-6.5 23</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24.5,-21.5,-5,-21.5</points>
<intersection>-24.5 2</intersection>
<intersection>-7 0</intersection>
<intersection>-5 25</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-24.5,-21.5,-24.5,0.5</points>
<intersection>-21.5 1</intersection>
<intersection>-16.5 12</intersection>
<intersection>-11.5 13</intersection>
<intersection>-6.5 14</intersection>
<intersection>-1.5 15</intersection>
<intersection>0.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-27,0.5,-24.5,0.5</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<intersection>-24.5 2</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-7,-24,-2.5,-24</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>-7 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-24.5,-16.5,-22,-16.5</points>
<intersection>-24.5 2</intersection>
<intersection>-22 19</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-24.5,-11.5,-22,-11.5</points>
<intersection>-24.5 2</intersection>
<intersection>-22 18</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-24.5,-6.5,-22,-6.5</points>
<intersection>-24.5 2</intersection>
<intersection>-22 17</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-24.5,-1.5,-22,-1.5</points>
<intersection>-24.5 2</intersection>
<intersection>-22 16</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-22,-2,-22,-1.5</points>
<connection>
<GID>26</GID>
<name>ENABLE_0</name></connection>
<intersection>-1.5 15</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>-22,-7,-22,-6.5</points>
<connection>
<GID>31</GID>
<name>ENABLE_0</name></connection>
<intersection>-6.5 14</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>-22,-12,-22,-11.5</points>
<connection>
<GID>34</GID>
<name>ENABLE_0</name></connection>
<intersection>-11.5 13</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>-22,-17,-22,-16.5</points>
<connection>
<GID>37</GID>
<name>ENABLE_0</name></connection>
<intersection>-16.5 12</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-7,-26,-6.5,-26</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>-7 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-7,-16.5,-5,-16.5</points>
<intersection>-7 0</intersection>
<intersection>-5 26</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-7,-6.5,-5,-6.5</points>
<intersection>-7 0</intersection>
<intersection>-5 28</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>-7,-11.5,-5,-11.5</points>
<intersection>-7 0</intersection>
<intersection>-5 27</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>-5,-21.5,-5,-21</points>
<connection>
<GID>38</GID>
<name>ENABLE_0</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>-5,-16.5,-5,-16</points>
<connection>
<GID>35</GID>
<name>ENABLE_0</name></connection>
<intersection>-16.5 22</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>-5,-11.5,-5,-11</points>
<connection>
<GID>32</GID>
<name>ENABLE_0</name></connection>
<intersection>-11.5 24</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>-5,-6.5,-5,-6</points>
<connection>
<GID>28</GID>
<name>ENABLE_0</name></connection>
<intersection>-6.5 23</intersection></vsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27,7.5,-26,7.5</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<connection>
<GID>55</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27,4,-26,4</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>-2.5,-26,-1.5,-26</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<connection>
<GID>61</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1019</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-4,-0.5,-4</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<connection>
<GID>1297</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1020</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-9,-0.5,-9</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<connection>
<GID>1298</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1021</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-14,-0.5,-14</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<connection>
<GID>1299</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1022</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-19,-0.5,-19</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<connection>
<GID>1300</GID>
<name>IN_0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-103.599,37.3091,207.518,-141.02</PageViewport>
<gate>
<ID>1</ID>
<type>BE_DECODER_3x8</type>
<position>-30,-28</position>
<input>
<ID>ENABLE</ID>46 </input>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>48 </input>
<input>
<ID>IN_2</ID>47 </input>
<output>
<ID>OUT_0</ID>102 </output>
<output>
<ID>OUT_1</ID>87 </output>
<output>
<ID>OUT_4</ID>86 </output>
<output>
<ID>OUT_5</ID>85 </output>
<output>
<ID>OUT_6</ID>84 </output>
<output>
<ID>OUT_7</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>4</ID>
<type>DA_FROM</type>
<position>-86.5,-6.5</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Cin  A</lparam></gate>
<gate>
<ID>27</ID>
<type>DA_FROM</type>
<position>-86.5,-8.5</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Data  C'</lparam></gate>
<gate>
<ID>30</ID>
<type>DA_FROM</type>
<position>-86.5,-11.5</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Cin  A</lparam></gate>
<gate>
<ID>33</ID>
<type>DA_FROM</type>
<position>-86.5,-13.5</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Self  B</lparam></gate>
<gate>
<ID>36</ID>
<type>DA_FROM</type>
<position>-86.5,-16.5</position>
<input>
<ID>IN_0</ID>34 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Self  B</lparam></gate>
<gate>
<ID>39</ID>
<type>DA_FROM</type>
<position>-86.5,-18.5</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Data  C'</lparam></gate>
<gate>
<ID>42</ID>
<type>EE_VDD</type>
<position>-34,-22.5</position>
<output>
<ID>OUT_0</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_AND2</type>
<position>-80.5,-7.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_AND2</type>
<position>-80.5,-12.5</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_AND2</type>
<position>-80.5,-17.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>58</ID>
<type>DA_FROM</type>
<position>-36,-28.5</position>
<input>
<ID>IN_0</ID>47 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>64</ID>
<type>AE_OR3</type>
<position>-73,-12.5</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>35 </input>
<input>
<ID>IN_2</ID>40 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>66</ID>
<type>DA_FROM</type>
<position>-36,-30.5</position>
<input>
<ID>IN_0</ID>48 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>70</ID>
<type>DE_TO</type>
<position>-67,-12.5</position>
<input>
<ID>IN_0</ID>45 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Cout</lparam></gate>
<gate>
<ID>71</ID>
<type>DA_FROM</type>
<position>-54,-6.5</position>
<input>
<ID>IN_0</ID>63 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Cin A</lparam></gate>
<gate>
<ID>76</ID>
<type>DA_FROM</type>
<position>-54,-8.5</position>
<input>
<ID>IN_0</ID>64 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C'</lparam></gate>
<gate>
<ID>80</ID>
<type>DA_FROM</type>
<position>-54,-11.5</position>
<input>
<ID>IN_0</ID>65 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>82</ID>
<type>DA_FROM</type>
<position>-54,-13.5</position>
<input>
<ID>IN_0</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>84</ID>
<type>DA_FROM</type>
<position>-54,-16.5</position>
<input>
<ID>IN_0</ID>68 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>86</ID>
<type>DA_FROM</type>
<position>-54,-18.5</position>
<input>
<ID>IN_0</ID>67 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C'</lparam></gate>
<gate>
<ID>88</ID>
<type>DA_FROM</type>
<position>-36,-32.5</position>
<input>
<ID>IN_0</ID>51 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>-52,-3</position>
<gparam>LABEL_TEXT Used NAND-NANDX</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>DE_TO</type>
<position>-5,-28.5</position>
<input>
<ID>IN_0</ID>61 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Mux 1</lparam></gate>
<gate>
<ID>102</ID>
<type>AA_LABEL</type>
<position>-102,10.5</position>
<gparam>LABEL_TEXT Key:</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>103</ID>
<type>DE_TO</type>
<position>-34.5,-12.5</position>
<input>
<ID>IN_0</ID>62 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Cout</lparam></gate>
<gate>
<ID>107</ID>
<type>DE_OR8</type>
<position>-12,-28.5</position>
<input>
<ID>IN_0</ID>83 </input>
<input>
<ID>IN_1</ID>84 </input>
<input>
<ID>IN_2</ID>85 </input>
<input>
<ID>IN_3</ID>86 </input>
<input>
<ID>IN_4</ID>103 </input>
<input>
<ID>IN_5</ID>103 </input>
<input>
<ID>IN_6</ID>102 </input>
<input>
<ID>IN_7</ID>87 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>108</ID>
<type>BI_NANDX3</type>
<position>-40.5,-12.5</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>70 </input>
<input>
<ID>IN_2</ID>71 </input>
<output>
<ID>OUT</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>109</ID>
<type>AA_LABEL</type>
<position>-102,7</position>
<gparam>LABEL_TEXT A = Cin</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>BA_NAND2</type>
<position>-48,-7.5</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>69 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>112</ID>
<type>BA_NAND2</type>
<position>-48,-12.5</position>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>BA_NAND2</type>
<position>-48,-17.5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>67 </input>
<output>
<ID>OUT</ID>71 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>114</ID>
<type>DA_FROM</type>
<position>-95.5,-27</position>
<input>
<ID>IN_0</ID>73 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>115</ID>
<type>DA_FROM</type>
<position>-95.5,-29</position>
<input>
<ID>IN_0</ID>72 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B'</lparam></gate>
<gate>
<ID>116</ID>
<type>FF_GND</type>
<position>-15,-34</position>
<output>
<ID>OUT_0</ID>103 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>117</ID>
<type>AE_OR2</type>
<position>-89.5,-28</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>72 </input>
<output>
<ID>OUT</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>118</ID>
<type>DE_TO</type>
<position>-83.5,-28</position>
<input>
<ID>IN_0</ID>74 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Mux 1</lparam></gate>
<gate>
<ID>119</ID>
<type>BE_DECODER_3x8</type>
<position>-22,-42.5</position>
<input>
<ID>ENABLE</ID>104 </input>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>106 </input>
<input>
<ID>IN_2</ID>105 </input>
<output>
<ID>OUT_2</ID>118 </output>
<output>
<ID>OUT_4</ID>117 </output>
<output>
<ID>OUT_5</ID>116 </output>
<output>
<ID>OUT_6</ID>115 </output>
<output>
<ID>OUT_7</ID>114 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>120</ID>
<type>BI_NANDX2</type>
<position>-57,-28</position>
<input>
<ID>IN_0</ID>75 </input>
<input>
<ID>IN_1</ID>76 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>121</ID>
<type>DA_FROM</type>
<position>-63,-27</position>
<input>
<ID>IN_0</ID>75 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A'</lparam></gate>
<gate>
<ID>122</ID>
<type>DA_FROM</type>
<position>-63,-29</position>
<input>
<ID>IN_0</ID>76 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>123</ID>
<type>DE_TO</type>
<position>-51,-28</position>
<input>
<ID>IN_0</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Mux 1</lparam></gate>
<gate>
<ID>124</ID>
<type>DA_FROM</type>
<position>-94.5,-41</position>
<input>
<ID>IN_0</ID>78 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>125</ID>
<type>DA_FROM</type>
<position>-94.5,-43</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C'</lparam></gate>
<gate>
<ID>126</ID>
<type>EE_VDD</type>
<position>-26,-37</position>
<output>
<ID>OUT_0</ID>104 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>127</ID>
<type>AA_AND2</type>
<position>-88.5,-42</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>128</ID>
<type>DA_FROM</type>
<position>-28,-43</position>
<input>
<ID>IN_0</ID>105 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>129</ID>
<type>AE_OR2</type>
<position>-81.5,-43</position>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>130</ID>
<type>DA_FROM</type>
<position>-87,-46</position>
<input>
<ID>IN_0</ID>81 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>131</ID>
<type>DE_TO</type>
<position>-75.5,-43</position>
<input>
<ID>IN_0</ID>82 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Mux 0</lparam></gate>
<gate>
<ID>132</ID>
<type>DA_FROM</type>
<position>-62,-41</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>133</ID>
<type>DA_FROM</type>
<position>-62,-43</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C'</lparam></gate>
<gate>
<ID>134</ID>
<type>DA_FROM</type>
<position>-28,-45</position>
<input>
<ID>IN_0</ID>106 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>135</ID>
<type>DA_FROM</type>
<position>-28,-47</position>
<input>
<ID>IN_0</ID>107 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>136</ID>
<type>DA_FROM</type>
<position>-54.5,-46</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>137</ID>
<type>DE_TO</type>
<position>-42,-43</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Mux 0</lparam></gate>
<gate>
<ID>138</ID>
<type>AA_LABEL</type>
<position>-102,4</position>
<gparam>LABEL_TEXT B = Self</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>139</ID>
<type>BA_NAND2</type>
<position>-56,-42</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT</ID>92 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>140</ID>
<type>DE_TO</type>
<position>-3.5,-42.5</position>
<input>
<ID>IN_0</ID>113 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Mux 0</lparam></gate>
<gate>
<ID>141</ID>
<type>BI_NANDX2</type>
<position>-48,-43</position>
<input>
<ID>IN_0</ID>92 </input>
<input>
<ID>IN_1</ID>91 </input>
<output>
<ID>OUT</ID>90 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>142</ID>
<type>AA_LABEL</type>
<position>-102,1</position>
<gparam>LABEL_TEXT C = Data</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>143</ID>
<type>BE_DECODER_3x8</type>
<position>-19,-13</position>
<input>
<ID>ENABLE</ID>93 </input>
<input>
<ID>IN_0</ID>96 </input>
<input>
<ID>IN_1</ID>95 </input>
<input>
<ID>IN_2</ID>94 </input>
<output>
<ID>OUT_2</ID>101 </output>
<output>
<ID>OUT_4</ID>100 </output>
<output>
<ID>OUT_6</ID>99 </output>
<output>
<ID>OUT_7</ID>98 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>144</ID>
<type>DE_OR8</type>
<position>-10.5,-42.5</position>
<input>
<ID>IN_0</ID>114 </input>
<input>
<ID>IN_1</ID>115 </input>
<input>
<ID>IN_2</ID>116 </input>
<input>
<ID>IN_3</ID>117 </input>
<input>
<ID>IN_4</ID>119 </input>
<input>
<ID>IN_5</ID>119 </input>
<input>
<ID>IN_6</ID>119 </input>
<input>
<ID>IN_7</ID>118 </input>
<output>
<ID>OUT</ID>113 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>145</ID>
<type>EE_VDD</type>
<position>-23,-7.5</position>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>146</ID>
<type>DA_FROM</type>
<position>-25,-13.5</position>
<input>
<ID>IN_0</ID>94 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>147</ID>
<type>DA_FROM</type>
<position>-25,-15.5</position>
<input>
<ID>IN_0</ID>95 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>148</ID>
<type>DA_FROM</type>
<position>-25,-17.5</position>
<input>
<ID>IN_0</ID>96 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>150</ID>
<type>AE_OR4</type>
<position>-7.5,-12.5</position>
<input>
<ID>IN_0</ID>98 </input>
<input>
<ID>IN_1</ID>99 </input>
<input>
<ID>IN_2</ID>100 </input>
<input>
<ID>IN_3</ID>101 </input>
<output>
<ID>OUT</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>151</ID>
<type>DE_TO</type>
<position>-0.5,-12.5</position>
<input>
<ID>IN_0</ID>97 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Cout</lparam></gate>
<gate>
<ID>152</ID>
<type>FF_GND</type>
<position>-13.5,-48</position>
<output>
<ID>OUT_0</ID>119 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_LABEL</type>
<position>-82.5,1</position>
<gparam>LABEL_TEXT Compare Logic</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-84.5,-6.5,-83.5,-6.5</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<connection>
<GID>4</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-84.5,-8.5,-83.5,-8.5</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<connection>
<GID>27</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-84.5,-13.5,-83.5,-13.5</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<connection>
<GID>33</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-84.5,-11.5,-83.5,-11.5</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<connection>
<GID>30</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-84.5,-18.5,-83.5,-18.5</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<connection>
<GID>39</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-84.5,-16.5,-83.5,-16.5</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<connection>
<GID>36</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-77.5,-12.5,-76,-12.5</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<connection>
<GID>64</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-76.5,-10.5,-76.5,-7.5</points>
<intersection>-10.5 1</intersection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-76.5,-10.5,-76,-10.5</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>-76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-77.5,-7.5,-76.5,-7.5</points>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<intersection>-76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-76.5,-17.5,-76.5,-14.5</points>
<intersection>-17.5 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-76.5,-14.5,-76,-14.5</points>
<connection>
<GID>64</GID>
<name>IN_2</name></connection>
<intersection>-76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-77.5,-17.5,-76.5,-17.5</points>
<connection>
<GID>56</GID>
<name>OUT</name></connection>
<intersection>-76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-70,-12.5,-69,-12.5</points>
<connection>
<GID>64</GID>
<name>OUT</name></connection>
<connection>
<GID>70</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-24.5,-34,-23.5</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34,-24.5,-33,-24.5</points>
<connection>
<GID>1</GID>
<name>ENABLE</name></connection>
<intersection>-34 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-34,-28.5,-33,-28.5</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>-33 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-33,-29.5,-33,-28.5</points>
<connection>
<GID>1</GID>
<name>IN_2</name></connection>
<intersection>-28.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-34,-30.5,-33,-30.5</points>
<connection>
<GID>1</GID>
<name>IN_1</name></connection>
<connection>
<GID>66</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33,-32.5,-33,-31.5</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34,-32.5,-33,-32.5</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>-33 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-8,-28.5,-7,-28.5</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<connection>
<GID>107</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-37.5,-12.5,-36.5,-12.5</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<connection>
<GID>108</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-52,-6.5,-51,-6.5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<connection>
<GID>71</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-52,-8.5,-51,-8.5</points>
<connection>
<GID>111</GID>
<name>IN_1</name></connection>
<connection>
<GID>76</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-52,-11.5,-51,-11.5</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<connection>
<GID>112</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-52,-13.5,-51,-13.5</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<connection>
<GID>112</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-52,-18.5,-51,-18.5</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<connection>
<GID>113</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-52,-16.5,-51,-16.5</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<connection>
<GID>113</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44,-10.5,-44,-7.5</points>
<intersection>-10.5 1</intersection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-44,-10.5,-43.5,-10.5</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>-44 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-45,-7.5,-44,-7.5</points>
<connection>
<GID>111</GID>
<name>OUT</name></connection>
<intersection>-44 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-45,-12.5,-43.5,-12.5</points>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<connection>
<GID>112</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44,-17.5,-44,-14.5</points>
<intersection>-17.5 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-44,-14.5,-43.5,-14.5</points>
<connection>
<GID>108</GID>
<name>IN_2</name></connection>
<intersection>-44 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-45,-17.5,-44,-17.5</points>
<connection>
<GID>113</GID>
<name>OUT</name></connection>
<intersection>-44 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-93.5,-29,-92.5,-29</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<connection>
<GID>117</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-93.5,-27,-92.5,-27</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<connection>
<GID>117</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-86.5,-28,-85.5,-28</points>
<connection>
<GID>117</GID>
<name>OUT</name></connection>
<connection>
<GID>118</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-61,-27,-60,-27</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<connection>
<GID>121</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-61,-29,-60,-29</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<connection>
<GID>122</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-54,-28,-53,-28</points>
<connection>
<GID>120</GID>
<name>OUT</name></connection>
<connection>
<GID>123</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-92.5,-41,-91.5,-41</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<connection>
<GID>127</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-92.5,-43,-91.5,-43</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<connection>
<GID>127</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-85.5,-42,-84.5,-42</points>
<connection>
<GID>127</GID>
<name>OUT</name></connection>
<connection>
<GID>129</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-84.5,-46,-84.5,-44</points>
<connection>
<GID>129</GID>
<name>IN_1</name></connection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-85,-46,-84.5,-46</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>-84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-78.5,-43,-77.5,-43</points>
<connection>
<GID>129</GID>
<name>OUT</name></connection>
<connection>
<GID>131</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-21,-25,-21,-24.5</points>
<intersection>-25 1</intersection>
<intersection>-24.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-21,-25,-15,-25</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>-21 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-27,-24.5,-21,-24.5</points>
<connection>
<GID>1</GID>
<name>OUT_7</name></connection>
<intersection>-21 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-21,-26,-21,-25.5</points>
<intersection>-26 1</intersection>
<intersection>-25.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-21,-26,-15,-26</points>
<connection>
<GID>107</GID>
<name>IN_1</name></connection>
<intersection>-21 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-27,-25.5,-21,-25.5</points>
<connection>
<GID>1</GID>
<name>OUT_6</name></connection>
<intersection>-21 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-21,-27,-21,-26.5</points>
<intersection>-27 1</intersection>
<intersection>-26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-21,-27,-15,-27</points>
<connection>
<GID>107</GID>
<name>IN_2</name></connection>
<intersection>-21 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-27,-26.5,-21,-26.5</points>
<connection>
<GID>1</GID>
<name>OUT_5</name></connection>
<intersection>-21 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-21,-28,-21,-27.5</points>
<intersection>-28 1</intersection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-21,-28,-15,-28</points>
<connection>
<GID>107</GID>
<name>IN_3</name></connection>
<intersection>-21 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-27,-27.5,-21,-27.5</points>
<connection>
<GID>1</GID>
<name>OUT_4</name></connection>
<intersection>-21 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-21,-30.5,-21,-29</points>
<intersection>-30.5 2</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-21,-29,-15,-29</points>
<connection>
<GID>107</GID>
<name>IN_7</name></connection>
<intersection>-21 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-27,-30.5,-21,-30.5</points>
<connection>
<GID>1</GID>
<name>OUT_1</name></connection>
<intersection>-21 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-60,-41,-59,-41</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<connection>
<GID>139</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-60,-43,-59,-43</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<connection>
<GID>139</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-45,-43,-44,-43</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<connection>
<GID>141</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52,-46,-52,-44</points>
<intersection>-46 1</intersection>
<intersection>-44 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-52.5,-46,-52,-46</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>-52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-52,-44,-51,-44</points>
<connection>
<GID>141</GID>
<name>IN_1</name></connection>
<intersection>-52 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<hsegment>
<ID>9</ID>
<points>-53,-42,-51,-42</points>
<connection>
<GID>139</GID>
<name>OUT</name></connection>
<connection>
<GID>141</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,-9.5,-23,-8.5</points>
<connection>
<GID>145</GID>
<name>OUT_0</name></connection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-23,-9.5,-22,-9.5</points>
<connection>
<GID>143</GID>
<name>ENABLE</name></connection>
<intersection>-23 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-23,-13.5,-22,-13.5</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>-22 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-22,-14.5,-22,-13.5</points>
<connection>
<GID>143</GID>
<name>IN_2</name></connection>
<intersection>-13.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-23,-15.5,-22,-15.5</points>
<connection>
<GID>143</GID>
<name>IN_1</name></connection>
<connection>
<GID>147</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22,-17.5,-22,-16.5</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-23,-17.5,-22,-17.5</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>-22 0</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<hsegment>
<ID>11</ID>
<points>-3.5,-12.5,-2.5,-12.5</points>
<connection>
<GID>150</GID>
<name>OUT</name></connection>
<connection>
<GID>151</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-16,-9.5,-10.5,-9.5</points>
<connection>
<GID>143</GID>
<name>OUT_7</name></connection>
<connection>
<GID>150</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-11.5,-10.5,-11.5</points>
<connection>
<GID>150</GID>
<name>IN_1</name></connection>
<intersection>-11.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-11.5,-11.5,-11.5,-10.5</points>
<intersection>-11.5 1</intersection>
<intersection>-10.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-16,-10.5,-11.5,-10.5</points>
<connection>
<GID>143</GID>
<name>OUT_6</name></connection>
<intersection>-11.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-13.5,-10.5,-13.5</points>
<connection>
<GID>150</GID>
<name>IN_2</name></connection>
<intersection>-11.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-11.5,-13.5,-11.5,-12.5</points>
<intersection>-13.5 1</intersection>
<intersection>-12.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-16,-12.5,-11.5,-12.5</points>
<connection>
<GID>143</GID>
<name>OUT_4</name></connection>
<intersection>-11.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-15.5,-10.5,-15.5</points>
<connection>
<GID>150</GID>
<name>IN_3</name></connection>
<intersection>-11.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-11.5,-15.5,-11.5,-14.5</points>
<intersection>-15.5 1</intersection>
<intersection>-14.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-16,-14.5,-11.5,-14.5</points>
<connection>
<GID>143</GID>
<name>OUT_2</name></connection>
<intersection>-11.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20.5,-31.5,-20.5,-30</points>
<intersection>-31.5 2</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-20.5,-30,-15,-30</points>
<connection>
<GID>107</GID>
<name>IN_6</name></connection>
<intersection>-20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-27,-31.5,-20.5,-31.5</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>-20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15,-33,-15,-31</points>
<connection>
<GID>107</GID>
<name>IN_4</name></connection>
<connection>
<GID>107</GID>
<name>IN_5</name></connection>
<connection>
<GID>116</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26,-39,-26,-38</points>
<connection>
<GID>126</GID>
<name>OUT_0</name></connection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-26,-39,-25,-39</points>
<connection>
<GID>119</GID>
<name>ENABLE</name></connection>
<intersection>-26 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-26,-43,-25,-43</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>-25 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-25,-44,-25,-43</points>
<connection>
<GID>119</GID>
<name>IN_2</name></connection>
<intersection>-43 1</intersection></vsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-26,-45,-25,-45</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<connection>
<GID>134</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25,-47,-25,-46</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>-47 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-26,-47,-25,-47</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>-25 0</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6.5,-42.5,-5.5,-42.5</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<connection>
<GID>144</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-19,-39,-13.5,-39</points>
<connection>
<GID>119</GID>
<name>OUT_7</name></connection>
<connection>
<GID>144</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-19,-40,-13.5,-40</points>
<connection>
<GID>119</GID>
<name>OUT_6</name></connection>
<connection>
<GID>144</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-19,-41,-13.5,-41</points>
<connection>
<GID>119</GID>
<name>OUT_5</name></connection>
<connection>
<GID>144</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-19,-42,-13.5,-42</points>
<connection>
<GID>119</GID>
<name>OUT_4</name></connection>
<connection>
<GID>144</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,-44,-16,-43</points>
<intersection>-44 2</intersection>
<intersection>-43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16,-43,-13.5,-43</points>
<connection>
<GID>144</GID>
<name>IN_7</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-19,-44,-16,-44</points>
<connection>
<GID>119</GID>
<name>OUT_2</name></connection>
<intersection>-16 0</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,-47,-13.5,-44</points>
<connection>
<GID>144</GID>
<name>IN_4</name></connection>
<connection>
<GID>144</GID>
<name>IN_5</name></connection>
<connection>
<GID>144</GID>
<name>IN_6</name></connection>
<connection>
<GID>152</GID>
<name>OUT_0</name></connection></vsegment></shape></wire></page 1>
<page 2>
<PageViewport>-51.7953,-3.694,119.319,-101.775</PageViewport>
<gate>
<ID>965</ID>
<type>BI_NANDX2</type>
<position>-20,-80.5</position>
<input>
<ID>IN_0</ID>741 </input>
<input>
<ID>IN_1</ID>740 </input>
<output>
<ID>OUT</ID>739 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>193</ID>
<type>HA_JUNC_2</type>
<position>76,-100.5</position>
<input>
<ID>N_in1</ID>153 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>966</ID>
<type>AE_SMALL_INVERTER</type>
<position>-27,-76.5</position>
<input>
<ID>IN_0</ID>735 </input>
<output>
<ID>OUT_0</ID>741 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>194</ID>
<type>HA_JUNC_2</type>
<position>76,-68</position>
<input>
<ID>N_in0</ID>167 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>195</ID>
<type>HA_JUNC_2</type>
<position>72.5,-71</position>
<input>
<ID>N_in0</ID>170 </input>
<input>
<ID>N_in1</ID>156 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>19.5,-12</position>
<gparam>LABEL_TEXT Used</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>582</ID>
<type>AA_LABEL</type>
<position>-31.5,-5</position>
<gparam>LABEL_TEXT Decision Logic</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>196</ID>
<type>HA_JUNC_2</type>
<position>72.5,-70</position>
<input>
<ID>N_in0</ID>169 </input>
<input>
<ID>N_in1</ID>157 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>197</ID>
<type>BA_NAND2</type>
<position>89,-87.5</position>
<input>
<ID>IN_0</ID>165 </input>
<input>
<ID>IN_1</ID>164 </input>
<output>
<ID>OUT</ID>160 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>HA_JUNC_2</type>
<position>69.5,-36.5</position>
<input>
<ID>N_in0</ID>495 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>198</ID>
<type>BA_NAND2</type>
<position>89,-92</position>
<input>
<ID>IN_0</ID>153 </input>
<input>
<ID>IN_1</ID>164 </input>
<output>
<ID>OUT</ID>161 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>585</ID>
<type>AA_LABEL</type>
<position>38.5,-14</position>
<gparam>LABEL_TEXT Mux0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>199</ID>
<type>HA_JUNC_2</type>
<position>99,-71</position>
<input>
<ID>N_in0</ID>156 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>200</ID>
<type>HA_JUNC_2</type>
<position>99,-70</position>
<input>
<ID>N_in0</ID>157 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>201</ID>
<type>BA_NAND2</type>
<position>89,-96.5</position>
<input>
<ID>IN_0</ID>165 </input>
<input>
<ID>IN_1</ID>153 </input>
<output>
<ID>OUT</ID>162 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>202</ID>
<type>DA_FROM</type>
<position>84.5,-82.5</position>
<input>
<ID>IN_0</ID>158 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>203</ID>
<type>BI_NANDX3</type>
<position>81.5,-92</position>
<input>
<ID>IN_0</ID>162 </input>
<input>
<ID>IN_1</ID>161 </input>
<input>
<ID>IN_2</ID>160 </input>
<output>
<ID>OUT</ID>163 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>204</ID>
<type>DA_FROM</type>
<position>84.5,-84.5</position>
<input>
<ID>IN_0</ID>159 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Reset</lparam></gate>
<gate>
<ID>205</ID>
<type>HA_JUNC_2</type>
<position>72.5,-92</position>
<input>
<ID>N_in0</ID>168 </input>
<input>
<ID>N_in1</ID>163 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>206</ID>
<type>AE_SMALL_INVERTER</type>
<position>97.5,-94.5</position>
<input>
<ID>IN_0</ID>155 </input>
<output>
<ID>OUT_0</ID>165 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>208</ID>
<type>HA_JUNC_2</type>
<position>101,-68</position>
<input>
<ID>N_in0</ID>173 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>210</ID>
<type>HE_JUNC_4</type>
<position>101,-92</position>
<input>
<ID>N_in0</ID>172 </input>
<input>
<ID>N_in2</ID>174 </input>
<input>
<ID>N_in3</ID>173 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>790</ID>
<type>AA_LABEL</type>
<position>72,-36.5</position>
<gparam>LABEL_TEXT Cin</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>212</ID>
<type>HA_JUNC_2</type>
<position>101,-100.5</position>
<input>
<ID>N_in1</ID>174 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>25</ID>
<type>HA_JUNC_2</type>
<position>13.5,-92</position>
<input>
<ID>N_in0</ID>56 </input>
<input>
<ID>N_in1</ID>134 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>606</ID>
<type>AA_LABEL</type>
<position>38.5,-15.5</position>
<gparam>LABEL_TEXT Mux1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AE_DFF_LOW</type>
<position>5.5,-79.5</position>
<input>
<ID>IN_0</ID>41 </input>
<output>
<ID>OUT_0</ID>39 </output>
<input>
<ID>clear</ID>50 </input>
<input>
<ID>clock</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>611</ID>
<type>AA_LABEL</type>
<position>45,-49.5</position>
<gparam>LABEL_TEXT Below</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>40</ID>
<type>DE_TO</type>
<position>5,-73</position>
<input>
<ID>IN_0</ID>39 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID N.3</lparam></gate>
<gate>
<ID>623</ID>
<type>AA_LABEL</type>
<position>46.5,-48.5</position>
<gparam>LABEL_TEXT Self</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>48</ID>
<type>AE_MUX_4x1</type>
<position>-2.5,-77.5</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>42 </input>
<input>
<ID>IN_2</ID>59 </input>
<input>
<ID>IN_3</ID>58 </input>
<output>
<ID>OUT</ID>41 </output>
<input>
<ID>SEL_0</ID>44 </input>
<input>
<ID>SEL_1</ID>43 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>52</ID>
<type>HA_JUNC_2</type>
<position>-10.5,-68</position>
<input>
<ID>N_in0</ID>39 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>632</ID>
<type>AA_LABEL</type>
<position>48,-49</position>
<gparam>LABEL_TEXT Data</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>637</ID>
<type>AE_OR2</type>
<position>-15.5,-28.5</position>
<input>
<ID>IN_0</ID>498 </input>
<input>
<ID>IN_1</ID>499 </input>
<output>
<ID>OUT</ID>502 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>60</ID>
<type>HA_JUNC_2</type>
<position>-10.5,-100.5</position>
<input>
<ID>N_in1</ID>58 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>62</ID>
<type>HA_JUNC_2</type>
<position>-8.5,-100.5</position>
<input>
<ID>N_in1</ID>42 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>646</ID>
<type>AA_LABEL</type>
<position>-8,-17.5</position>
<gparam>LABEL_TEXT Mux0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>HA_JUNC_2</type>
<position>-8.5,-68</position>
<input>
<ID>N_in0</ID>42 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>649</ID>
<type>AE_OR2</type>
<position>-15.5,-23.5</position>
<input>
<ID>IN_0</ID>497 </input>
<input>
<ID>IN_1</ID>498 </input>
<output>
<ID>OUT</ID>501 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>72</ID>
<type>HA_JUNC_2</type>
<position>-9.5,-100.5</position>
<input>
<ID>N_in1</ID>39 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>73</ID>
<type>HA_JUNC_2</type>
<position>-9.5,-68</position>
<input>
<ID>N_in0</ID>59 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>74</ID>
<type>HA_JUNC_2</type>
<position>-13,-71</position>
<input>
<ID>N_in0</ID>109 </input>
<input>
<ID>N_in1</ID>43 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>HA_JUNC_2</type>
<position>-13,-70</position>
<input>
<ID>N_in0</ID>108 </input>
<input>
<ID>N_in1</ID>44 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>656</ID>
<type>AA_LABEL</type>
<position>-8,-19</position>
<gparam>LABEL_TEXT Mux1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>BA_NAND2</type>
<position>3.5,-87.5</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>56 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>78</ID>
<type>BA_NAND2</type>
<position>3.5,-92</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>56 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>79</ID>
<type>HA_JUNC_2</type>
<position>13.5,-71</position>
<input>
<ID>N_in0</ID>43 </input>
<input>
<ID>N_in1</ID>133 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>HA_JUNC_2</type>
<position>13.5,-70</position>
<input>
<ID>N_in0</ID>44 </input>
<input>
<ID>N_in1</ID>132 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>661</ID>
<type>AI_XOR2</type>
<position>-21.5,-21</position>
<input>
<ID>IN_0</ID>503 </input>
<input>
<ID>IN_1</ID>500 </input>
<output>
<ID>OUT</ID>497 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>83</ID>
<type>BA_NAND2</type>
<position>3.5,-96.5</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>663</ID>
<type>AE_DFF_LOW</type>
<position>61.5,-24</position>
<input>
<ID>IN_0</ID>485 </input>
<output>
<ID>OUT_0</ID>484 </output>
<input>
<ID>clear</ID>490 </input>
<input>
<ID>clock</ID>489 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>85</ID>
<type>DA_FROM</type>
<position>-1,-82.5</position>
<input>
<ID>IN_0</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>665</ID>
<type>AA_LABEL</type>
<position>-8,-40</position>
<gparam>LABEL_TEXT Cout Final</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>BI_NANDX3</type>
<position>-4,-92</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>53 </input>
<input>
<ID>IN_2</ID>52 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>667</ID>
<type>DE_TO</type>
<position>61,-17.5</position>
<input>
<ID>IN_0</ID>484 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID N.n</lparam></gate>
<gate>
<ID>89</ID>
<type>DA_FROM</type>
<position>-1,-84.5</position>
<input>
<ID>IN_0</ID>50 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Reset</lparam></gate>
<gate>
<ID>670</ID>
<type>AE_MUX_4x1</type>
<position>53.5,-22</position>
<input>
<ID>IN_0</ID>484 </input>
<input>
<ID>IN_1</ID>486 </input>
<input>
<ID>IN_2</ID>505 </input>
<input>
<ID>IN_3</ID>504 </input>
<output>
<ID>OUT</ID>485 </output>
<input>
<ID>SEL_0</ID>488 </input>
<input>
<ID>SEL_1</ID>487 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>91</ID>
<type>HA_JUNC_2</type>
<position>-13,-92</position>
<input>
<ID>N_in0</ID>60 </input>
<input>
<ID>N_in1</ID>55 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>672</ID>
<type>AA_LABEL</type>
<position>-33.5,-61.5</position>
<gparam>LABEL_TEXT 4-Bit Unit</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>93</ID>
<type>AE_SMALL_INVERTER</type>
<position>12,-94.5</position>
<input>
<ID>IN_0</ID>42 </input>
<output>
<ID>OUT_0</ID>57 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>94</ID>
<type>HA_JUNC_2</type>
<position>42,-92</position>
<input>
<ID>N_in0</ID>128 </input>
<input>
<ID>N_in1</ID>150 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>674</ID>
<type>HA_JUNC_2</type>
<position>45.5,-12.5</position>
<input>
<ID>N_in0</ID>484 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>95</ID>
<type>AE_DFF_LOW</type>
<position>34,-79.5</position>
<input>
<ID>IN_0</ID>111 </input>
<output>
<ID>OUT_0</ID>110 </output>
<input>
<ID>clear</ID>123 </input>
<input>
<ID>clock</ID>122 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>96</ID>
<type>DE_TO</type>
<position>33.5,-73</position>
<input>
<ID>IN_0</ID>110 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID N.2</lparam></gate>
<gate>
<ID>97</ID>
<type>AE_MUX_4x1</type>
<position>26,-77.5</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>112 </input>
<input>
<ID>IN_2</ID>131 </input>
<input>
<ID>IN_3</ID>130 </input>
<output>
<ID>OUT</ID>111 </output>
<input>
<ID>SEL_0</ID>121 </input>
<input>
<ID>SEL_1</ID>120 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>677</ID>
<type>HA_JUNC_2</type>
<position>45.5,-45</position>
<input>
<ID>N_in1</ID>504 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>98</ID>
<type>HA_JUNC_2</type>
<position>18,-68</position>
<input>
<ID>N_in0</ID>110 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>99</ID>
<type>HA_JUNC_2</type>
<position>18,-100.5</position>
<input>
<ID>N_in1</ID>130 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>100</ID>
<type>HA_JUNC_2</type>
<position>20,-100.5</position>
<input>
<ID>N_in1</ID>112 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>680</ID>
<type>HA_JUNC_2</type>
<position>47.5,-45</position>
<input>
<ID>N_in1</ID>486 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>101</ID>
<type>HA_JUNC_2</type>
<position>20,-68</position>
<input>
<ID>N_in0</ID>112 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>683</ID>
<type>HA_JUNC_2</type>
<position>47.5,-12.5</position>
<input>
<ID>N_in0</ID>486 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>104</ID>
<type>HA_JUNC_2</type>
<position>19,-100.5</position>
<input>
<ID>N_in1</ID>110 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>105</ID>
<type>HA_JUNC_2</type>
<position>19,-68</position>
<input>
<ID>N_in0</ID>131 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>685</ID>
<type>HA_JUNC_2</type>
<position>46.5,-45</position>
<input>
<ID>N_in1</ID>484 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>106</ID>
<type>HA_JUNC_2</type>
<position>15.5,-71</position>
<input>
<ID>N_in0</ID>133 </input>
<input>
<ID>N_in1</ID>120 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>686</ID>
<type>HA_JUNC_2</type>
<position>46.5,-12.5</position>
<input>
<ID>N_in0</ID>505 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>687</ID>
<type>HA_JUNC_2</type>
<position>43,-15.5</position>
<input>
<ID>N_in1</ID>487 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>688</ID>
<type>HA_JUNC_2</type>
<position>43,-14.5</position>
<input>
<ID>N_in1</ID>488 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>689</ID>
<type>BA_NAND2</type>
<position>59.5,-32</position>
<input>
<ID>IN_0</ID>496 </input>
<input>
<ID>IN_1</ID>495 </input>
<output>
<ID>OUT</ID>491 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>110</ID>
<type>HA_JUNC_2</type>
<position>15.5,-70</position>
<input>
<ID>N_in0</ID>132 </input>
<input>
<ID>N_in1</ID>121 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>690</ID>
<type>BA_NAND2</type>
<position>59.5,-36.5</position>
<input>
<ID>IN_0</ID>484 </input>
<input>
<ID>IN_1</ID>495 </input>
<output>
<ID>OUT</ID>492 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>691</ID>
<type>HA_JUNC_2</type>
<position>69.5,-15.5</position>
<input>
<ID>N_in0</ID>487 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>692</ID>
<type>HA_JUNC_2</type>
<position>69.5,-14.5</position>
<input>
<ID>N_in0</ID>488 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>693</ID>
<type>BA_NAND2</type>
<position>59.5,-41</position>
<input>
<ID>IN_0</ID>496 </input>
<input>
<ID>IN_1</ID>484 </input>
<output>
<ID>OUT</ID>493 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>694</ID>
<type>DA_FROM</type>
<position>55,-27</position>
<input>
<ID>IN_0</ID>489 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>695</ID>
<type>BI_NANDX3</type>
<position>52,-36.5</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>492 </input>
<input>
<ID>IN_2</ID>491 </input>
<output>
<ID>OUT</ID>494 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>696</ID>
<type>DA_FROM</type>
<position>55,-29</position>
<input>
<ID>IN_0</ID>490 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Reset</lparam></gate>
<gate>
<ID>697</ID>
<type>HA_JUNC_2</type>
<position>43,-36.5</position>
<input>
<ID>N_in1</ID>494 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>698</ID>
<type>AA_LABEL</type>
<position>41.5,-5.5</position>
<gparam>LABEL_TEXT 1-Bit Cell</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>700</ID>
<type>AE_SMALL_INVERTER</type>
<position>68,-39</position>
<input>
<ID>IN_0</ID>486 </input>
<output>
<ID>OUT_0</ID>496 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>701</ID>
<type>AA_LABEL</type>
<position>39,-36.5</position>
<gparam>LABEL_TEXT Cout</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>714</ID>
<type>HA_JUNC_2</type>
<position>-25,-16</position>
<input>
<ID>N_in0</ID>503 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>715</ID>
<type>HA_JUNC_2</type>
<position>-25,-48.5</position>
<input>
<ID>N_in1</ID>500 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>716</ID>
<type>AE_SMALL_INVERTER</type>
<position>-22,-29.5</position>
<input>
<ID>IN_0</ID>503 </input>
<output>
<ID>OUT_0</ID>499 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>717</ID>
<type>HA_JUNC_2</type>
<position>-10.5,-18</position>
<input>
<ID>N_in0</ID>501 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>718</ID>
<type>HA_JUNC_2</type>
<position>-10.5,-19</position>
<input>
<ID>N_in0</ID>502 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>719</ID>
<type>HA_JUNC_2</type>
<position>-10.5,-40</position>
<input>
<ID>N_in0</ID>500 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>720</ID>
<type>HA_JUNC_2</type>
<position>-26,-16</position>
<input>
<ID>N_in0</ID>498 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>721</ID>
<type>HA_JUNC_2</type>
<position>-26,-48.5</position>
<input>
<ID>N_in1</ID>498 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>722</ID>
<type>AA_LABEL</type>
<position>46.5,-10</position>
<gparam>LABEL_TEXT Above</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>723</ID>
<type>AA_LABEL</type>
<position>45,-10</position>
<gparam>LABEL_TEXT Self</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>724</ID>
<type>AA_LABEL</type>
<position>48,-10</position>
<gparam>LABEL_TEXT Data</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>725</ID>
<type>AA_LABEL</type>
<position>-26,-52.5</position>
<gparam>LABEL_TEXT R/W</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>726</ID>
<type>AA_LABEL</type>
<position>-24.5,-51.5</position>
<gparam>LABEL_TEXT CF</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>727</ID>
<type>AA_LABEL</type>
<position>-26,-13.5</position>
<gparam>LABEL_TEXT R/W</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>728</ID>
<type>AA_LABEL</type>
<position>-24.5,-13.5</position>
<gparam>LABEL_TEXT Above CF</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>149</ID>
<type>BA_NAND2</type>
<position>32,-87.5</position>
<input>
<ID>IN_0</ID>129 </input>
<input>
<ID>IN_1</ID>128 </input>
<output>
<ID>OUT</ID>124 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>733</ID>
<type>AA_LABEL</type>
<position>27.5,-17.5</position>
<gparam>LABEL_TEXT Mux0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>154</ID>
<type>BA_NAND2</type>
<position>32,-92</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>128 </input>
<output>
<ID>OUT</ID>125 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>155</ID>
<type>HA_JUNC_2</type>
<position>42,-71</position>
<input>
<ID>N_in0</ID>120 </input>
<input>
<ID>N_in1</ID>152 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>735</ID>
<type>AA_LABEL</type>
<position>27.5,-19</position>
<gparam>LABEL_TEXT Mux1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>156</ID>
<type>HA_JUNC_2</type>
<position>42,-70</position>
<input>
<ID>N_in0</ID>121 </input>
<input>
<ID>N_in1</ID>151 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>BA_NAND2</type>
<position>32,-96.5</position>
<input>
<ID>IN_0</ID>129 </input>
<input>
<ID>IN_1</ID>110 </input>
<output>
<ID>OUT</ID>126 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>737</ID>
<type>AA_LABEL</type>
<position>27.5,-40</position>
<gparam>LABEL_TEXT Cout Final</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>158</ID>
<type>DA_FROM</type>
<position>27.5,-82.5</position>
<input>
<ID>IN_0</ID>122 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>738</ID>
<type>HA_JUNC_2</type>
<position>10.5,-16</position>
<input>
<ID>N_in0</ID>598 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>159</ID>
<type>BI_NANDX3</type>
<position>24.5,-92</position>
<input>
<ID>IN_0</ID>126 </input>
<input>
<ID>IN_1</ID>125 </input>
<input>
<ID>IN_2</ID>124 </input>
<output>
<ID>OUT</ID>127 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>739</ID>
<type>HA_JUNC_2</type>
<position>10.5,-48.5</position>
<input>
<ID>N_in1</ID>589 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>160</ID>
<type>DA_FROM</type>
<position>27.5,-84.5</position>
<input>
<ID>IN_0</ID>123 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Reset</lparam></gate>
<gate>
<ID>161</ID>
<type>HA_JUNC_2</type>
<position>15.5,-92</position>
<input>
<ID>N_in0</ID>134 </input>
<input>
<ID>N_in1</ID>127 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>741</ID>
<type>HA_JUNC_2</type>
<position>25,-18</position>
<input>
<ID>N_in0</ID>596 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>162</ID>
<type>AE_SMALL_INVERTER</type>
<position>40.5,-94.5</position>
<input>
<ID>IN_0</ID>112 </input>
<output>
<ID>OUT_0</ID>129 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>742</ID>
<type>HA_JUNC_2</type>
<position>25,-19</position>
<input>
<ID>N_in0</ID>597 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>163</ID>
<type>HA_JUNC_2</type>
<position>70.5,-92</position>
<input>
<ID>N_in0</ID>146 </input>
<input>
<ID>N_in1</ID>168 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>743</ID>
<type>HA_JUNC_2</type>
<position>25,-40</position>
<input>
<ID>N_in0</ID>589 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>164</ID>
<type>AE_DFF_LOW</type>
<position>62.5,-79.5</position>
<input>
<ID>IN_0</ID>136 </input>
<output>
<ID>OUT_0</ID>135 </output>
<input>
<ID>clear</ID>141 </input>
<input>
<ID>clock</ID>140 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>744</ID>
<type>HA_JUNC_2</type>
<position>9.5,-16</position>
<input>
<ID>N_in0</ID>587 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>165</ID>
<type>DE_TO</type>
<position>62,-73</position>
<input>
<ID>IN_0</ID>135 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID N.1</lparam></gate>
<gate>
<ID>745</ID>
<type>HA_JUNC_2</type>
<position>9.5,-48.5</position>
<input>
<ID>N_in1</ID>587 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>166</ID>
<type>AE_MUX_4x1</type>
<position>54.5,-77.5</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>137 </input>
<input>
<ID>IN_2</ID>149 </input>
<input>
<ID>IN_3</ID>148 </input>
<output>
<ID>OUT</ID>136 </output>
<input>
<ID>SEL_0</ID>139 </input>
<input>
<ID>SEL_1</ID>138 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>746</ID>
<type>AA_LABEL</type>
<position>9.5,-52.5</position>
<gparam>LABEL_TEXT R/W</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>167</ID>
<type>HA_JUNC_2</type>
<position>46.5,-68</position>
<input>
<ID>N_in0</ID>135 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>747</ID>
<type>AA_LABEL</type>
<position>11,-51.5</position>
<gparam>LABEL_TEXT CF</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>168</ID>
<type>HA_JUNC_2</type>
<position>46.5,-100.5</position>
<input>
<ID>N_in1</ID>148 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>748</ID>
<type>AA_LABEL</type>
<position>9.5,-13.5</position>
<gparam>LABEL_TEXT R/W</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>169</ID>
<type>HA_JUNC_2</type>
<position>48.5,-100.5</position>
<input>
<ID>N_in1</ID>137 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>749</ID>
<type>AA_LABEL</type>
<position>11,-13.5</position>
<gparam>LABEL_TEXT Above CF</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>170</ID>
<type>HA_JUNC_2</type>
<position>48.5,-68</position>
<input>
<ID>N_in0</ID>137 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>171</ID>
<type>HA_JUNC_2</type>
<position>47.5,-100.5</position>
<input>
<ID>N_in1</ID>135 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>751</ID>
<type>AO_XNOR2</type>
<position>14,-21</position>
<input>
<ID>IN_0</ID>598 </input>
<input>
<ID>IN_1</ID>589 </input>
<output>
<ID>OUT</ID>594 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>172</ID>
<type>HA_JUNC_2</type>
<position>47.5,-68</position>
<input>
<ID>N_in0</ID>149 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>173</ID>
<type>HA_JUNC_2</type>
<position>44,-71</position>
<input>
<ID>N_in0</ID>152 </input>
<input>
<ID>N_in1</ID>138 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>753</ID>
<type>BI_NANDX2</type>
<position>20,-23.5</position>
<input>
<ID>IN_0</ID>594 </input>
<input>
<ID>IN_1</ID>599 </input>
<output>
<ID>OUT</ID>596 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>174</ID>
<type>HA_JUNC_2</type>
<position>44,-70</position>
<input>
<ID>N_in0</ID>151 </input>
<input>
<ID>N_in1</ID>139 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>754</ID>
<type>BI_NANDX2</type>
<position>20,-28.5</position>
<input>
<ID>IN_0</ID>599 </input>
<input>
<ID>IN_1</ID>598 </input>
<output>
<ID>OUT</ID>597 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>175</ID>
<type>BA_NAND2</type>
<position>60.5,-87.5</position>
<input>
<ID>IN_0</ID>147 </input>
<input>
<ID>IN_1</ID>146 </input>
<output>
<ID>OUT</ID>142 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>176</ID>
<type>BA_NAND2</type>
<position>60.5,-92</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>146 </input>
<output>
<ID>OUT</ID>143 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>177</ID>
<type>HA_JUNC_2</type>
<position>70.5,-71</position>
<input>
<ID>N_in0</ID>138 </input>
<input>
<ID>N_in1</ID>170 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>757</ID>
<type>AE_SMALL_INVERTER</type>
<position>13,-24.5</position>
<input>
<ID>IN_0</ID>587 </input>
<output>
<ID>OUT_0</ID>599 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>178</ID>
<type>HA_JUNC_2</type>
<position>70.5,-70</position>
<input>
<ID>N_in0</ID>139 </input>
<input>
<ID>N_in1</ID>169 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>179</ID>
<type>BA_NAND2</type>
<position>60.5,-96.5</position>
<input>
<ID>IN_0</ID>147 </input>
<input>
<ID>IN_1</ID>135 </input>
<output>
<ID>OUT</ID>144 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>952</ID>
<type>HA_JUNC_2</type>
<position>-29.5,-68</position>
<input>
<ID>N_in0</ID>740 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>180</ID>
<type>DA_FROM</type>
<position>56,-82.5</position>
<input>
<ID>IN_0</ID>140 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>953</ID>
<type>HA_JUNC_2</type>
<position>-29.5,-100.5</position>
<input>
<ID>N_in1</ID>736 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>181</ID>
<type>BI_NANDX3</type>
<position>53,-92</position>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>143 </input>
<input>
<ID>IN_2</ID>142 </input>
<output>
<ID>OUT</ID>145 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>954</ID>
<type>HA_JUNC_2</type>
<position>-15,-70</position>
<input>
<ID>N_in0</ID>738 </input>
<input>
<ID>N_in1</ID>108 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>182</ID>
<type>DA_FROM</type>
<position>56,-84.5</position>
<input>
<ID>IN_0</ID>141 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Reset</lparam></gate>
<gate>
<ID>955</ID>
<type>HA_JUNC_2</type>
<position>-15,-71</position>
<input>
<ID>N_in0</ID>739 </input>
<input>
<ID>N_in1</ID>109 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>183</ID>
<type>HA_JUNC_2</type>
<position>44,-92</position>
<input>
<ID>N_in0</ID>150 </input>
<input>
<ID>N_in1</ID>145 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>956</ID>
<type>HA_JUNC_2</type>
<position>-15,-92</position>
<input>
<ID>N_in0</ID>736 </input>
<input>
<ID>N_in1</ID>60 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>184</ID>
<type>AE_SMALL_INVERTER</type>
<position>69,-94.5</position>
<input>
<ID>IN_0</ID>137 </input>
<output>
<ID>OUT_0</ID>147 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>957</ID>
<type>HA_JUNC_2</type>
<position>-30.5,-68</position>
<input>
<ID>N_in0</ID>735 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>185</ID>
<type>HA_JUNC_2</type>
<position>99,-92</position>
<input>
<ID>N_in0</ID>164 </input>
<input>
<ID>N_in1</ID>172 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>958</ID>
<type>HA_JUNC_2</type>
<position>-30.5,-100.5</position>
<input>
<ID>N_in1</ID>735 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>186</ID>
<type>AE_DFF_LOW</type>
<position>91,-79.5</position>
<input>
<ID>IN_0</ID>154 </input>
<output>
<ID>OUT_0</ID>153 </output>
<input>
<ID>clear</ID>159 </input>
<input>
<ID>clock</ID>158 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>187</ID>
<type>DE_TO</type>
<position>90.5,-73</position>
<input>
<ID>IN_0</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID N.0</lparam></gate>
<gate>
<ID>188</ID>
<type>AE_MUX_4x1</type>
<position>83,-77.5</position>
<input>
<ID>IN_0</ID>153 </input>
<input>
<ID>IN_1</ID>155 </input>
<input>
<ID>IN_2</ID>167 </input>
<input>
<ID>IN_3</ID>166 </input>
<output>
<ID>OUT</ID>154 </output>
<input>
<ID>SEL_0</ID>157 </input>
<input>
<ID>SEL_1</ID>156 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>189</ID>
<type>HA_JUNC_2</type>
<position>75,-68</position>
<input>
<ID>N_in0</ID>153 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>190</ID>
<type>HA_JUNC_2</type>
<position>75,-100.5</position>
<input>
<ID>N_in1</ID>166 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>963</ID>
<type>AO_XNOR2</type>
<position>-26,-73</position>
<input>
<ID>IN_0</ID>740 </input>
<input>
<ID>IN_1</ID>736 </input>
<output>
<ID>OUT</ID>737 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>191</ID>
<type>HA_JUNC_2</type>
<position>77,-100.5</position>
<input>
<ID>N_in1</ID>155 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>964</ID>
<type>BI_NANDX2</type>
<position>-20,-75.5</position>
<input>
<ID>IN_0</ID>737 </input>
<input>
<ID>IN_1</ID>741 </input>
<output>
<ID>OUT</ID>738 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>192</ID>
<type>HA_JUNC_2</type>
<position>77,-68</position>
<input>
<ID>N_in0</ID>155 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<wire>
<ID>587</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-47.5,9.5,-17</points>
<connection>
<GID>745</GID>
<name>N_in1</name></connection>
<connection>
<GID>744</GID>
<name>N_in0</name></connection>
<intersection>-24.5 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>9.5,-24.5,11,-24.5</points>
<connection>
<GID>757</GID>
<name>IN_0</name></connection>
<intersection>9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>589</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>10,-40,24,-40</points>
<connection>
<GID>743</GID>
<name>N_in0</name></connection>
<intersection>10 8</intersection>
<intersection>10.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>10.5,-47.5,10.5,-40</points>
<connection>
<GID>739</GID>
<name>N_in1</name></connection>
<intersection>-40 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>10,-40,10,-22</points>
<intersection>-40 2</intersection>
<intersection>-22 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>10,-22,11,-22</points>
<connection>
<GID>751</GID>
<name>IN_1</name></connection>
<intersection>10 8</intersection></hsegment></shape></wire>
<wire>
<ID>594</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-22.5,17,-21</points>
<connection>
<GID>753</GID>
<name>IN_0</name></connection>
<connection>
<GID>751</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>596</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-23.5,23,-18</points>
<connection>
<GID>753</GID>
<name>OUT</name></connection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-18,24,-18</points>
<connection>
<GID>741</GID>
<name>N_in0</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>597</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-28.5,24,-19</points>
<connection>
<GID>742</GID>
<name>N_in0</name></connection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>23,-28.5,24,-28.5</points>
<connection>
<GID>754</GID>
<name>OUT</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>598</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-29.5,10.5,-17</points>
<connection>
<GID>738</GID>
<name>N_in0</name></connection>
<intersection>-29.5 3</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10.5,-20,11,-20</points>
<connection>
<GID>751</GID>
<name>IN_0</name></connection>
<intersection>10.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>10.5,-29.5,17,-29.5</points>
<connection>
<GID>754</GID>
<name>IN_1</name></connection>
<intersection>10.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>599</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-24.5,17,-24.5</points>
<connection>
<GID>753</GID>
<name>IN_1</name></connection>
<connection>
<GID>757</GID>
<name>OUT_0</name></connection>
<intersection>16 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>16,-27.5,16,-24.5</points>
<intersection>-27.5 8</intersection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>16,-27.5,17,-27.5</points>
<connection>
<GID>754</GID>
<name>IN_0</name></connection>
<intersection>16 7</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-100,9.5,-75</points>
<intersection>-100 2</intersection>
<intersection>-95.5 14</intersection>
<intersection>-77.5 7</intersection>
<intersection>-75 30</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-10.5,-100,9.5,-100</points>
<intersection>-10.5 4</intersection>
<intersection>-9.5 17</intersection>
<intersection>9.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-10.5,-100,-10.5,-69</points>
<connection>
<GID>52</GID>
<name>N_in0</name></connection>
<intersection>-100 2</intersection>
<intersection>-80.5 9</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>8.5,-77.5,9.5,-77.5</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>9.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-10.5,-80.5,-5.5,-80.5</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>-10.5 4</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>6.5,-95.5,9.5,-95.5</points>
<connection>
<GID>83</GID>
<name>IN_1</name></connection>
<intersection>6.5 27</intersection>
<intersection>9.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>-9.5,-100,-9.5,-99.5</points>
<connection>
<GID>72</GID>
<name>N_in1</name></connection>
<intersection>-100 2</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>6.5,-95.5,6.5,-93</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>-95.5 14</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>3,-75,9.5,-75</points>
<intersection>3 32</intersection>
<intersection>9.5 0</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>3,-75,3,-73</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>-75 30</intersection></vsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0.5,-77.5,2.5,-77.5</points>
<connection>
<GID>48</GID>
<name>OUT</name></connection>
<connection>
<GID>29</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8.5,-100.5,-8.5,-69</points>
<connection>
<GID>62</GID>
<name>N_in1</name></connection>
<connection>
<GID>68</GID>
<name>N_in0</name></connection>
<intersection>-100.5 6</intersection>
<intersection>-78.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-8.5,-78.5,-5.5,-78.5</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>-8.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-8.5,-100.5,14,-100.5</points>
<intersection>-8.5 0</intersection>
<intersection>14 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>14,-100.5,14,-94.5</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>-100.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2.5,-72.5,-2.5,-71</points>
<connection>
<GID>48</GID>
<name>SEL_1</name></connection>
<intersection>-71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12,-71,12.5,-71</points>
<connection>
<GID>74</GID>
<name>N_in1</name></connection>
<connection>
<GID>79</GID>
<name>N_in0</name></connection>
<intersection>-2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1.5,-72.5,-1.5,-70</points>
<connection>
<GID>48</GID>
<name>SEL_0</name></connection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12,-70,12.5,-70</points>
<connection>
<GID>75</GID>
<name>N_in1</name></connection>
<connection>
<GID>81</GID>
<name>N_in0</name></connection>
<intersection>-1.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,-82.5,2.5,-80.5</points>
<connection>
<GID>29</GID>
<name>clock</name></connection>
<intersection>-82.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1,-82.5,2.5,-82.5</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,-84.5,5.5,-83.5</points>
<connection>
<GID>29</GID>
<name>clear</name></connection>
<intersection>-84.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>1,-84.5,5.5,-84.5</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-0.5,-90,-0.5,-87.5</points>
<intersection>-90 1</intersection>
<intersection>-87.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1,-90,-0.5,-90</points>
<connection>
<GID>87</GID>
<name>IN_2</name></connection>
<intersection>-0.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-0.5,-87.5,0.5,-87.5</points>
<connection>
<GID>77</GID>
<name>OUT</name></connection>
<intersection>-0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-92,0.5,-92</points>
<connection>
<GID>87</GID>
<name>IN_1</name></connection>
<connection>
<GID>78</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-0.5,-96.5,-0.5,-94</points>
<intersection>-96.5 1</intersection>
<intersection>-94 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-0.5,-96.5,0.5,-96.5</points>
<connection>
<GID>83</GID>
<name>OUT</name></connection>
<intersection>-0.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1,-94,-0.5,-94</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>-0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-12,-92,-7,-92</points>
<connection>
<GID>91</GID>
<name>N_in1</name></connection>
<connection>
<GID>87</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-92,10.5,-86.5</points>
<intersection>-92 8</intersection>
<intersection>-91 1</intersection>
<intersection>-86.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6.5,-91,10.5,-91</points>
<connection>
<GID>78</GID>
<name>IN_1</name></connection>
<intersection>10.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>6.5,-86.5,10.5,-86.5</points>
<connection>
<GID>77</GID>
<name>IN_1</name></connection>
<intersection>10.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>10.5,-92,12.5,-92</points>
<connection>
<GID>25</GID>
<name>N_in0</name></connection>
<intersection>10.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8.5,-97.5,8.5,-88.5</points>
<intersection>-97.5 3</intersection>
<intersection>-94.5 2</intersection>
<intersection>-88.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6.5,-88.5,8.5,-88.5</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-94.5,10,-94.5</points>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>6.5,-97.5,8.5,-97.5</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>8.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,-99.5,-11,-74.5</points>
<intersection>-99.5 2</intersection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-11,-74.5,-5.5,-74.5</points>
<connection>
<GID>48</GID>
<name>IN_3</name></connection>
<intersection>-11 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-11,-99.5,-10.5,-99.5</points>
<connection>
<GID>60</GID>
<name>N_in1</name></connection>
<intersection>-11 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9.5,-76.5,-9.5,-69</points>
<connection>
<GID>73</GID>
<name>N_in0</name></connection>
<intersection>-76.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-9.5,-76.5,-5.5,-76.5</points>
<connection>
<GID>48</GID>
<name>IN_2</name></connection>
<intersection>-9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,-92,-14,-92</points>
<connection>
<GID>91</GID>
<name>N_in0</name></connection>
<connection>
<GID>956</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>484</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-44.5,65.5,-19.5</points>
<intersection>-44.5 2</intersection>
<intersection>-40 14</intersection>
<intersection>-22 7</intersection>
<intersection>-19.5 30</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-44.5,65.5,-44.5</points>
<intersection>45.5 4</intersection>
<intersection>46.5 17</intersection>
<intersection>65.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>45.5,-44.5,45.5,-13.5</points>
<connection>
<GID>674</GID>
<name>N_in0</name></connection>
<intersection>-44.5 2</intersection>
<intersection>-25 9</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>64.5,-22,65.5,-22</points>
<connection>
<GID>663</GID>
<name>OUT_0</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>45.5,-25,50.5,-25</points>
<connection>
<GID>670</GID>
<name>IN_0</name></connection>
<intersection>45.5 4</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>62.5,-40,65.5,-40</points>
<connection>
<GID>693</GID>
<name>IN_1</name></connection>
<intersection>62.5 27</intersection>
<intersection>65.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>46.5,-44.5,46.5,-44</points>
<connection>
<GID>685</GID>
<name>N_in1</name></connection>
<intersection>-44.5 2</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>62.5,-40,62.5,-37.5</points>
<connection>
<GID>690</GID>
<name>IN_0</name></connection>
<intersection>-40 14</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>59,-19.5,65.5,-19.5</points>
<intersection>59 32</intersection>
<intersection>65.5 0</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>59,-19.5,59,-17.5</points>
<connection>
<GID>667</GID>
<name>IN_0</name></connection>
<intersection>-19.5 30</intersection></vsegment></shape></wire>
<wire>
<ID>485</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56.5,-22,58.5,-22</points>
<connection>
<GID>670</GID>
<name>OUT</name></connection>
<connection>
<GID>663</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>486</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-45,47.5,-13.5</points>
<connection>
<GID>680</GID>
<name>N_in1</name></connection>
<connection>
<GID>683</GID>
<name>N_in0</name></connection>
<intersection>-45 6</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>47.5,-23,50.5,-23</points>
<connection>
<GID>670</GID>
<name>IN_1</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>47.5,-45,70,-45</points>
<intersection>47.5 0</intersection>
<intersection>70 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>70,-45,70,-39</points>
<connection>
<GID>700</GID>
<name>IN_0</name></connection>
<intersection>-45 6</intersection></vsegment></shape></wire>
<wire>
<ID>487</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-17,53.5,-15.5</points>
<connection>
<GID>670</GID>
<name>SEL_1</name></connection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-15.5,68.5,-15.5</points>
<connection>
<GID>687</GID>
<name>N_in1</name></connection>
<connection>
<GID>691</GID>
<name>N_in0</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>488</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-17,54.5,-14.5</points>
<connection>
<GID>670</GID>
<name>SEL_0</name></connection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-14.5,68.5,-14.5</points>
<connection>
<GID>688</GID>
<name>N_in1</name></connection>
<connection>
<GID>692</GID>
<name>N_in0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>489</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-27,58.5,-25</points>
<connection>
<GID>663</GID>
<name>clock</name></connection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57,-27,58.5,-27</points>
<connection>
<GID>694</GID>
<name>IN_0</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>490</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-29,61.5,-28</points>
<connection>
<GID>663</GID>
<name>clear</name></connection>
<intersection>-29 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>57,-29,61.5,-29</points>
<connection>
<GID>696</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>491</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-34.5,55.5,-32</points>
<intersection>-34.5 1</intersection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-34.5,55.5,-34.5</points>
<connection>
<GID>695</GID>
<name>IN_2</name></connection>
<intersection>55.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55.5,-32,56.5,-32</points>
<connection>
<GID>689</GID>
<name>OUT</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>492</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-36.5,56.5,-36.5</points>
<connection>
<GID>695</GID>
<name>IN_1</name></connection>
<connection>
<GID>690</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>493</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-41,55.5,-38.5</points>
<intersection>-41 1</intersection>
<intersection>-38.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,-41,56.5,-41</points>
<connection>
<GID>693</GID>
<name>OUT</name></connection>
<intersection>55.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55,-38.5,55.5,-38.5</points>
<connection>
<GID>695</GID>
<name>IN_0</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>494</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>44,-36.5,49,-36.5</points>
<connection>
<GID>697</GID>
<name>N_in1</name></connection>
<connection>
<GID>695</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,-70,-14,-70</points>
<connection>
<GID>75</GID>
<name>N_in0</name></connection>
<connection>
<GID>954</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,-71,-14,-71</points>
<connection>
<GID>74</GID>
<name>N_in0</name></connection>
<connection>
<GID>955</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>495</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-36.5,66.5,-31</points>
<intersection>-36.5 8</intersection>
<intersection>-35.5 1</intersection>
<intersection>-31 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-35.5,66.5,-35.5</points>
<connection>
<GID>690</GID>
<name>IN_1</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>62.5,-31,66.5,-31</points>
<connection>
<GID>689</GID>
<name>IN_1</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>66.5,-36.5,68.5,-36.5</points>
<connection>
<GID>5</GID>
<name>N_in0</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>496</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-42,64.5,-33</points>
<intersection>-42 3</intersection>
<intersection>-39 2</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-33,64.5,-33</points>
<connection>
<GID>689</GID>
<name>IN_0</name></connection>
<intersection>64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-39,66,-39</points>
<connection>
<GID>700</GID>
<name>OUT_0</name></connection>
<intersection>64.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>62.5,-42,64.5,-42</points>
<connection>
<GID>693</GID>
<name>IN_0</name></connection>
<intersection>64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-100,38,-75</points>
<intersection>-100 2</intersection>
<intersection>-95.5 14</intersection>
<intersection>-77.5 7</intersection>
<intersection>-75 30</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>18,-100,38,-100</points>
<intersection>18 4</intersection>
<intersection>19 17</intersection>
<intersection>38 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>18,-100,18,-69</points>
<connection>
<GID>98</GID>
<name>N_in0</name></connection>
<intersection>-100 2</intersection>
<intersection>-80.5 9</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>37,-77.5,38,-77.5</points>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>18,-80.5,23,-80.5</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>18 4</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>35,-95.5,38,-95.5</points>
<connection>
<GID>157</GID>
<name>IN_1</name></connection>
<intersection>35 27</intersection>
<intersection>38 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>19,-100,19,-99.5</points>
<connection>
<GID>104</GID>
<name>N_in1</name></connection>
<intersection>-100 2</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>35,-95.5,35,-93</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>-95.5 14</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>31.5,-75,38,-75</points>
<intersection>31.5 32</intersection>
<intersection>38 0</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>31.5,-75,31.5,-73</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>-75 30</intersection></vsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,-77.5,31,-77.5</points>
<connection>
<GID>97</GID>
<name>OUT</name></connection>
<connection>
<GID>95</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>497</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-18.5,-22.5,-18.5,-21</points>
<connection>
<GID>661</GID>
<name>OUT</name></connection>
<connection>
<GID>649</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-100.5,20,-69</points>
<connection>
<GID>101</GID>
<name>N_in0</name></connection>
<connection>
<GID>100</GID>
<name>N_in1</name></connection>
<intersection>-100.5 6</intersection>
<intersection>-78.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>20,-78.5,23,-78.5</points>
<connection>
<GID>97</GID>
<name>IN_1</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>20,-100.5,42.5,-100.5</points>
<intersection>20 0</intersection>
<intersection>42.5 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>42.5,-100.5,42.5,-94.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>-100.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>498</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26,-47.5,-26,-17</points>
<connection>
<GID>721</GID>
<name>N_in1</name></connection>
<connection>
<GID>720</GID>
<name>N_in0</name></connection>
<intersection>-27.5 3</intersection>
<intersection>-24.5 15</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-26,-27.5,-18.5,-27.5</points>
<connection>
<GID>637</GID>
<name>IN_0</name></connection>
<intersection>-26 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-26,-24.5,-18.5,-24.5</points>
<connection>
<GID>649</GID>
<name>IN_1</name></connection>
<intersection>-26 0</intersection></hsegment></shape></wire>
<wire>
<ID>499</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-20,-29.5,-18.5,-29.5</points>
<connection>
<GID>637</GID>
<name>IN_1</name></connection>
<connection>
<GID>716</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>500</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25.5,-40,-25.5,-22</points>
<intersection>-40 2</intersection>
<intersection>-22 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-25.5,-40,-11.5,-40</points>
<connection>
<GID>719</GID>
<name>N_in0</name></connection>
<intersection>-25.5 0</intersection>
<intersection>-25 7</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-25.5,-22,-24.5,-22</points>
<connection>
<GID>661</GID>
<name>IN_1</name></connection>
<intersection>-25.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-25,-47.5,-25,-40</points>
<connection>
<GID>715</GID>
<name>N_in1</name></connection>
<intersection>-40 2</intersection></vsegment></shape></wire>
<wire>
<ID>501</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12.5,-23.5,-12.5,-18</points>
<connection>
<GID>649</GID>
<name>OUT</name></connection>
<intersection>-18 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-12.5,-18,-11.5,-18</points>
<connection>
<GID>717</GID>
<name>N_in0</name></connection>
<intersection>-12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>502</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11.5,-28.5,-11.5,-19</points>
<connection>
<GID>718</GID>
<name>N_in0</name></connection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12.5,-28.5,-11.5,-28.5</points>
<connection>
<GID>637</GID>
<name>OUT</name></connection>
<intersection>-11.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>503</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25,-29.5,-25,-17</points>
<connection>
<GID>714</GID>
<name>N_in0</name></connection>
<intersection>-29.5 4</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25,-20,-24.5,-20</points>
<connection>
<GID>661</GID>
<name>IN_0</name></connection>
<intersection>-25 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-25,-29.5,-24,-29.5</points>
<connection>
<GID>716</GID>
<name>IN_0</name></connection>
<intersection>-25 0</intersection></hsegment></shape></wire>
<wire>
<ID>504</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-44,45,-19</points>
<intersection>-44 2</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-19,50.5,-19</points>
<connection>
<GID>670</GID>
<name>IN_3</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-44,45.5,-44</points>
<connection>
<GID>677</GID>
<name>N_in1</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>505</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-21,46.5,-13.5</points>
<connection>
<GID>686</GID>
<name>N_in0</name></connection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-21,50.5,-21</points>
<connection>
<GID>670</GID>
<name>IN_2</name></connection>
<intersection>46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-72.5,26,-71</points>
<connection>
<GID>97</GID>
<name>SEL_1</name></connection>
<intersection>-71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16.5,-71,41,-71</points>
<connection>
<GID>155</GID>
<name>N_in0</name></connection>
<connection>
<GID>106</GID>
<name>N_in1</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-72.5,27,-70</points>
<connection>
<GID>97</GID>
<name>SEL_0</name></connection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16.5,-70,41,-70</points>
<connection>
<GID>156</GID>
<name>N_in0</name></connection>
<connection>
<GID>110</GID>
<name>N_in1</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-82.5,31,-80.5</points>
<connection>
<GID>95</GID>
<name>clock</name></connection>
<intersection>-82.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-82.5,31,-82.5</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-84.5,34,-83.5</points>
<connection>
<GID>95</GID>
<name>clear</name></connection>
<intersection>-84.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-84.5,34,-84.5</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-90,28,-87.5</points>
<intersection>-90 1</intersection>
<intersection>-87.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-90,28,-90</points>
<connection>
<GID>159</GID>
<name>IN_2</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28,-87.5,29,-87.5</points>
<connection>
<GID>149</GID>
<name>OUT</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-92,29,-92</points>
<connection>
<GID>159</GID>
<name>IN_1</name></connection>
<connection>
<GID>154</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-96.5,28,-94</points>
<intersection>-96.5 1</intersection>
<intersection>-94 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-96.5,29,-96.5</points>
<connection>
<GID>157</GID>
<name>OUT</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-94,28,-94</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>16.5,-92,21.5,-92</points>
<connection>
<GID>161</GID>
<name>N_in1</name></connection>
<connection>
<GID>159</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-92,39,-86.5</points>
<intersection>-92 8</intersection>
<intersection>-91 1</intersection>
<intersection>-86.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-91,39,-91</points>
<connection>
<GID>154</GID>
<name>IN_1</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>35,-86.5,39,-86.5</points>
<connection>
<GID>149</GID>
<name>IN_1</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>39,-92,41,-92</points>
<connection>
<GID>94</GID>
<name>N_in0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-97.5,37,-88.5</points>
<intersection>-97.5 3</intersection>
<intersection>-94.5 2</intersection>
<intersection>-88.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-88.5,37,-88.5</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37,-94.5,38.5,-94.5</points>
<connection>
<GID>162</GID>
<name>OUT_0</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>35,-97.5,37,-97.5</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-99.5,17.5,-74.5</points>
<intersection>-99.5 2</intersection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-74.5,23,-74.5</points>
<connection>
<GID>97</GID>
<name>IN_3</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-99.5,18,-99.5</points>
<connection>
<GID>99</GID>
<name>N_in1</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-76.5,19,-69</points>
<connection>
<GID>105</GID>
<name>N_in0</name></connection>
<intersection>-76.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-76.5,23,-76.5</points>
<connection>
<GID>97</GID>
<name>IN_2</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-70,14.5,-70</points>
<connection>
<GID>81</GID>
<name>N_in1</name></connection>
<connection>
<GID>110</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-71,14.5,-71</points>
<connection>
<GID>79</GID>
<name>N_in1</name></connection>
<connection>
<GID>106</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-92,14.5,-92</points>
<connection>
<GID>25</GID>
<name>N_in1</name></connection>
<connection>
<GID>161</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-100,66.5,-75</points>
<intersection>-100 2</intersection>
<intersection>-95.5 14</intersection>
<intersection>-77.5 7</intersection>
<intersection>-75 30</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>46.5,-100,66.5,-100</points>
<intersection>46.5 4</intersection>
<intersection>47.5 17</intersection>
<intersection>66.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>46.5,-100,46.5,-69</points>
<connection>
<GID>167</GID>
<name>N_in0</name></connection>
<intersection>-100 2</intersection>
<intersection>-80.5 9</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>65.5,-77.5,66.5,-77.5</points>
<connection>
<GID>164</GID>
<name>OUT_0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>46.5,-80.5,51.5,-80.5</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>46.5 4</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>63.5,-95.5,66.5,-95.5</points>
<connection>
<GID>179</GID>
<name>IN_1</name></connection>
<intersection>63.5 27</intersection>
<intersection>66.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>47.5,-100,47.5,-99.5</points>
<connection>
<GID>171</GID>
<name>N_in1</name></connection>
<intersection>-100 2</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>63.5,-95.5,63.5,-93</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>-95.5 14</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>60,-75,66.5,-75</points>
<intersection>60 32</intersection>
<intersection>66.5 0</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>60,-75,60,-73</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>-75 30</intersection></vsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57.5,-77.5,59.5,-77.5</points>
<connection>
<GID>166</GID>
<name>OUT</name></connection>
<connection>
<GID>164</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,-100.5,48.5,-69</points>
<connection>
<GID>170</GID>
<name>N_in0</name></connection>
<connection>
<GID>169</GID>
<name>N_in1</name></connection>
<intersection>-100.5 6</intersection>
<intersection>-78.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-78.5,51.5,-78.5</points>
<connection>
<GID>166</GID>
<name>IN_1</name></connection>
<intersection>48.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>48.5,-100.5,71,-100.5</points>
<intersection>48.5 0</intersection>
<intersection>71 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>71,-100.5,71,-94.5</points>
<connection>
<GID>184</GID>
<name>IN_0</name></connection>
<intersection>-100.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-72.5,54.5,-71</points>
<connection>
<GID>166</GID>
<name>SEL_1</name></connection>
<intersection>-71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-71,69.5,-71</points>
<connection>
<GID>177</GID>
<name>N_in0</name></connection>
<connection>
<GID>173</GID>
<name>N_in1</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-72.5,55.5,-70</points>
<connection>
<GID>166</GID>
<name>SEL_0</name></connection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-70,69.5,-70</points>
<connection>
<GID>178</GID>
<name>N_in0</name></connection>
<connection>
<GID>174</GID>
<name>N_in1</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-82.5,59.5,-80.5</points>
<connection>
<GID>164</GID>
<name>clock</name></connection>
<intersection>-82.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,-82.5,59.5,-82.5</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-84.5,62.5,-83.5</points>
<connection>
<GID>164</GID>
<name>clear</name></connection>
<intersection>-84.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>58,-84.5,62.5,-84.5</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-90,56.5,-87.5</points>
<intersection>-90 1</intersection>
<intersection>-87.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-90,56.5,-90</points>
<connection>
<GID>181</GID>
<name>IN_2</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-87.5,57.5,-87.5</points>
<connection>
<GID>175</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56,-92,57.5,-92</points>
<connection>
<GID>181</GID>
<name>IN_1</name></connection>
<connection>
<GID>176</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-96.5,56.5,-94</points>
<intersection>-96.5 1</intersection>
<intersection>-94 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,-96.5,57.5,-96.5</points>
<connection>
<GID>179</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-94,56.5,-94</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>45,-92,50,-92</points>
<connection>
<GID>183</GID>
<name>N_in1</name></connection>
<connection>
<GID>181</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-92,67.5,-86.5</points>
<intersection>-92 8</intersection>
<intersection>-91 1</intersection>
<intersection>-86.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-91,67.5,-91</points>
<connection>
<GID>176</GID>
<name>IN_1</name></connection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>63.5,-86.5,67.5,-86.5</points>
<connection>
<GID>175</GID>
<name>IN_1</name></connection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>67.5,-92,69.5,-92</points>
<connection>
<GID>163</GID>
<name>N_in0</name></connection>
<intersection>67.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-97.5,65.5,-88.5</points>
<intersection>-97.5 3</intersection>
<intersection>-94.5 2</intersection>
<intersection>-88.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-88.5,65.5,-88.5</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65.5,-94.5,67,-94.5</points>
<connection>
<GID>184</GID>
<name>OUT_0</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>63.5,-97.5,65.5,-97.5</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-99.5,46,-74.5</points>
<intersection>-99.5 2</intersection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-74.5,51.5,-74.5</points>
<connection>
<GID>166</GID>
<name>IN_3</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46,-99.5,46.5,-99.5</points>
<connection>
<GID>168</GID>
<name>N_in1</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-76.5,47.5,-69</points>
<connection>
<GID>172</GID>
<name>N_in0</name></connection>
<intersection>-76.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-76.5,51.5,-76.5</points>
<connection>
<GID>166</GID>
<name>IN_2</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-92,43,-92</points>
<connection>
<GID>94</GID>
<name>N_in1</name></connection>
<connection>
<GID>183</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-70,43,-70</points>
<connection>
<GID>156</GID>
<name>N_in1</name></connection>
<connection>
<GID>174</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-71,43,-71</points>
<connection>
<GID>155</GID>
<name>N_in1</name></connection>
<connection>
<GID>173</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-100,95,-75</points>
<intersection>-100 2</intersection>
<intersection>-95.5 14</intersection>
<intersection>-77.5 7</intersection>
<intersection>-75 30</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>75,-100,95,-100</points>
<intersection>75 4</intersection>
<intersection>76 17</intersection>
<intersection>95 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>75,-100,75,-69</points>
<connection>
<GID>189</GID>
<name>N_in0</name></connection>
<intersection>-100 2</intersection>
<intersection>-80.5 9</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>94,-77.5,95,-77.5</points>
<connection>
<GID>186</GID>
<name>OUT_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>75,-80.5,80,-80.5</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>75 4</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>92,-95.5,95,-95.5</points>
<connection>
<GID>201</GID>
<name>IN_1</name></connection>
<intersection>92 27</intersection>
<intersection>95 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>76,-100,76,-99.5</points>
<connection>
<GID>193</GID>
<name>N_in1</name></connection>
<intersection>-100 2</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>92,-95.5,92,-93</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>-95.5 14</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>88.5,-75,95,-75</points>
<intersection>88.5 32</intersection>
<intersection>95 0</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>88.5,-75,88.5,-73</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>-75 30</intersection></vsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86,-77.5,88,-77.5</points>
<connection>
<GID>188</GID>
<name>OUT</name></connection>
<connection>
<GID>186</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-100.5,77,-69</points>
<connection>
<GID>192</GID>
<name>N_in0</name></connection>
<connection>
<GID>191</GID>
<name>N_in1</name></connection>
<intersection>-100.5 6</intersection>
<intersection>-78.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>77,-78.5,80,-78.5</points>
<connection>
<GID>188</GID>
<name>IN_1</name></connection>
<intersection>77 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>77,-100.5,99.5,-100.5</points>
<intersection>77 0</intersection>
<intersection>99.5 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>99.5,-100.5,99.5,-94.5</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>-100.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-72.5,83,-71</points>
<connection>
<GID>188</GID>
<name>SEL_1</name></connection>
<intersection>-71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-71,98,-71</points>
<connection>
<GID>199</GID>
<name>N_in0</name></connection>
<connection>
<GID>195</GID>
<name>N_in1</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>735</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30.5,-99.5,-30.5,-69</points>
<connection>
<GID>958</GID>
<name>N_in1</name></connection>
<connection>
<GID>957</GID>
<name>N_in0</name></connection>
<intersection>-76.5 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>-30.5,-76.5,-29,-76.5</points>
<connection>
<GID>966</GID>
<name>IN_0</name></connection>
<intersection>-30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>736</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-30,-92,-16,-92</points>
<connection>
<GID>956</GID>
<name>N_in0</name></connection>
<intersection>-30 8</intersection>
<intersection>-29.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-29.5,-99.5,-29.5,-92</points>
<connection>
<GID>953</GID>
<name>N_in1</name></connection>
<intersection>-92 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-30,-92,-30,-74</points>
<intersection>-92 2</intersection>
<intersection>-74 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-30,-74,-29,-74</points>
<connection>
<GID>963</GID>
<name>IN_1</name></connection>
<intersection>-30 8</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-72.5,84,-70</points>
<connection>
<GID>188</GID>
<name>SEL_0</name></connection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-70,98,-70</points>
<connection>
<GID>200</GID>
<name>N_in0</name></connection>
<connection>
<GID>196</GID>
<name>N_in1</name></connection>
<intersection>84 0</intersection></hsegment></shape></wire>
<wire>
<ID>737</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,-74.5,-23,-73</points>
<connection>
<GID>964</GID>
<name>IN_0</name></connection>
<connection>
<GID>963</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-82.5,88,-80.5</points>
<connection>
<GID>186</GID>
<name>clock</name></connection>
<intersection>-82.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86.5,-82.5,88,-82.5</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>88 0</intersection></hsegment></shape></wire>
<wire>
<ID>738</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-17,-75.5,-17,-70</points>
<connection>
<GID>964</GID>
<name>OUT</name></connection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-17,-70,-16,-70</points>
<connection>
<GID>954</GID>
<name>N_in0</name></connection>
<intersection>-17 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-84.5,91,-83.5</points>
<connection>
<GID>186</GID>
<name>clear</name></connection>
<intersection>-84.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-84.5,91,-84.5</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<intersection>91 0</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-90,85,-87.5</points>
<intersection>-90 1</intersection>
<intersection>-87.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84.5,-90,85,-90</points>
<connection>
<GID>203</GID>
<name>IN_2</name></connection>
<intersection>85 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>85,-87.5,86,-87.5</points>
<connection>
<GID>197</GID>
<name>OUT</name></connection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>739</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,-80.5,-16,-71</points>
<connection>
<GID>955</GID>
<name>N_in0</name></connection>
<intersection>-80.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-17,-80.5,-16,-80.5</points>
<connection>
<GID>965</GID>
<name>OUT</name></connection>
<intersection>-16 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,-92,86,-92</points>
<connection>
<GID>203</GID>
<name>IN_1</name></connection>
<connection>
<GID>198</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>740</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29.5,-81.5,-29.5,-69</points>
<connection>
<GID>952</GID>
<name>N_in0</name></connection>
<intersection>-81.5 3</intersection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29.5,-72,-29,-72</points>
<connection>
<GID>963</GID>
<name>IN_0</name></connection>
<intersection>-29.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-29.5,-81.5,-23,-81.5</points>
<connection>
<GID>965</GID>
<name>IN_1</name></connection>
<intersection>-29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-96.5,85,-94</points>
<intersection>-96.5 1</intersection>
<intersection>-94 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-96.5,86,-96.5</points>
<connection>
<GID>201</GID>
<name>OUT</name></connection>
<intersection>85 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84.5,-94,85,-94</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>741</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-25,-76.5,-23,-76.5</points>
<connection>
<GID>966</GID>
<name>OUT_0</name></connection>
<connection>
<GID>964</GID>
<name>IN_1</name></connection>
<intersection>-24 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-24,-79.5,-24,-76.5</points>
<intersection>-79.5 8</intersection>
<intersection>-76.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-24,-79.5,-23,-79.5</points>
<connection>
<GID>965</GID>
<name>IN_0</name></connection>
<intersection>-24 7</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>73.5,-92,78.5,-92</points>
<connection>
<GID>205</GID>
<name>N_in1</name></connection>
<connection>
<GID>203</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96,-92,96,-86.5</points>
<intersection>-92 8</intersection>
<intersection>-91 1</intersection>
<intersection>-86.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92,-91,96,-91</points>
<connection>
<GID>198</GID>
<name>IN_1</name></connection>
<intersection>96 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>92,-86.5,96,-86.5</points>
<connection>
<GID>197</GID>
<name>IN_1</name></connection>
<intersection>96 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>96,-92,98,-92</points>
<connection>
<GID>185</GID>
<name>N_in0</name></connection>
<intersection>96 0</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94,-97.5,94,-88.5</points>
<intersection>-97.5 3</intersection>
<intersection>-94.5 2</intersection>
<intersection>-88.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92,-88.5,94,-88.5</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>94 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94,-94.5,95.5,-94.5</points>
<connection>
<GID>206</GID>
<name>OUT_0</name></connection>
<intersection>94 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>92,-97.5,94,-97.5</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<intersection>94 0</intersection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-99.5,74.5,-74.5</points>
<intersection>-99.5 2</intersection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-74.5,80,-74.5</points>
<connection>
<GID>188</GID>
<name>IN_3</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74.5,-99.5,75,-99.5</points>
<connection>
<GID>190</GID>
<name>N_in1</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-76.5,76,-69</points>
<connection>
<GID>194</GID>
<name>N_in0</name></connection>
<intersection>-76.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-76.5,80,-76.5</points>
<connection>
<GID>188</GID>
<name>IN_2</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,-92,71.5,-92</points>
<connection>
<GID>205</GID>
<name>N_in0</name></connection>
<connection>
<GID>163</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,-70,71.5,-70</points>
<connection>
<GID>196</GID>
<name>N_in0</name></connection>
<connection>
<GID>178</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,-71,71.5,-71</points>
<connection>
<GID>195</GID>
<name>N_in0</name></connection>
<connection>
<GID>177</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-92,100,-92</points>
<connection>
<GID>210</GID>
<name>N_in0</name></connection>
<connection>
<GID>185</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-91,101,-69</points>
<connection>
<GID>210</GID>
<name>N_in3</name></connection>
<connection>
<GID>208</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-99.5,101,-93</points>
<connection>
<GID>210</GID>
<name>N_in2</name></connection>
<connection>
<GID>212</GID>
<name>N_in1</name></connection></vsegment></shape></wire></page 2>
<page 3>
<PageViewport>6.14136,252.151,796.49,-200.868</PageViewport>
<gate>
<ID>213</ID>
<type>HA_JUNC_2</type>
<position>186.5,148</position>
<input>
<ID>N_in0</ID>346 </input>
<input>
<ID>N_in1</ID>230 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>214</ID>
<type>BI_NANDX2</type>
<position>90.5,168</position>
<input>
<ID>IN_0</ID>257 </input>
<input>
<ID>IN_1</ID>256 </input>
<output>
<ID>OUT</ID>255 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>215</ID>
<type>HA_JUNC_2</type>
<position>186.5,180.5</position>
<input>
<ID>N_in0</ID>244 </input>
<input>
<ID>N_in1</ID>574 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>216</ID>
<type>AE_SMALL_INVERTER</type>
<position>83.5,172</position>
<input>
<ID>IN_0</ID>251 </input>
<output>
<ID>OUT_0</ID>257 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>217</ID>
<type>HA_JUNC_2</type>
<position>183,177.5</position>
<input>
<ID>N_in0</ID>247 </input>
<input>
<ID>N_in1</ID>233 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>218</ID>
<type>HA_JUNC_2</type>
<position>183,178.5</position>
<input>
<ID>N_in0</ID>246 </input>
<input>
<ID>N_in1</ID>234 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>219</ID>
<type>BA_NAND2</type>
<position>199.5,161</position>
<input>
<ID>IN_0</ID>242 </input>
<input>
<ID>IN_1</ID>241 </input>
<output>
<ID>OUT</ID>237 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>220</ID>
<type>BA_NAND2</type>
<position>199.5,156.5</position>
<input>
<ID>IN_0</ID>230 </input>
<input>
<ID>IN_1</ID>241 </input>
<output>
<ID>OUT</ID>238 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>221</ID>
<type>HA_JUNC_2</type>
<position>209.5,177.5</position>
<input>
<ID>N_in0</ID>233 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>222</ID>
<type>HA_JUNC_2</type>
<position>209.5,178.5</position>
<input>
<ID>N_in0</ID>234 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>223</ID>
<type>BA_NAND2</type>
<position>199.5,152</position>
<input>
<ID>IN_0</ID>242 </input>
<input>
<ID>IN_1</ID>230 </input>
<output>
<ID>OUT</ID>239 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>224</ID>
<type>DA_FROM</type>
<position>195,166</position>
<input>
<ID>IN_0</ID>235 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>225</ID>
<type>BI_NANDX3</type>
<position>192,156.5</position>
<input>
<ID>IN_0</ID>239 </input>
<input>
<ID>IN_1</ID>238 </input>
<input>
<ID>IN_2</ID>237 </input>
<output>
<ID>OUT</ID>240 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>226</ID>
<type>DA_FROM</type>
<position>195,164</position>
<input>
<ID>IN_0</ID>236 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Reset</lparam></gate>
<gate>
<ID>227</ID>
<type>HA_JUNC_2</type>
<position>183,156.5</position>
<input>
<ID>N_in0</ID>245 </input>
<input>
<ID>N_in1</ID>240 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>228</ID>
<type>AE_SMALL_INVERTER</type>
<position>208,154</position>
<input>
<ID>IN_0</ID>232 </input>
<output>
<ID>OUT_0</ID>242 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>229</ID>
<type>HA_JUNC_2</type>
<position>211.5,180.5</position>
<input>
<ID>N_in0</ID>249 </input>
<input>
<ID>N_in1</ID>574 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>230</ID>
<type>HE_JUNC_4</type>
<position>211.5,156.5</position>
<input>
<ID>N_in0</ID>248 </input>
<input>
<ID>N_in2</ID>250 </input>
<input>
<ID>N_in3</ID>249 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>231</ID>
<type>HA_JUNC_2</type>
<position>211.5,148</position>
<input>
<ID>N_in0</ID>345 </input>
<input>
<ID>N_in1</ID>250 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>232</ID>
<type>HA_JUNC_2</type>
<position>124,156.5</position>
<input>
<ID>N_in0</ID>187 </input>
<input>
<ID>N_in1</ID>211 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>233</ID>
<type>AE_DFF_LOW</type>
<position>116,169</position>
<input>
<ID>IN_0</ID>177 </input>
<output>
<ID>OUT_0</ID>176 </output>
<input>
<ID>clear</ID>182 </input>
<input>
<ID>clock</ID>181 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>234</ID>
<type>DE_TO</type>
<position>115.5,175.5</position>
<input>
<ID>IN_0</ID>176 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 0.3</lparam></gate>
<gate>
<ID>235</ID>
<type>AE_MUX_4x1</type>
<position>108,171</position>
<input>
<ID>IN_0</ID>176 </input>
<input>
<ID>IN_1</ID>178 </input>
<input>
<ID>IN_2</ID>190 </input>
<input>
<ID>IN_3</ID>189 </input>
<output>
<ID>OUT</ID>177 </output>
<input>
<ID>SEL_0</ID>180 </input>
<input>
<ID>SEL_1</ID>179 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>236</ID>
<type>HA_JUNC_2</type>
<position>100,180.5</position>
<input>
<ID>N_in0</ID>176 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>237</ID>
<type>HA_JUNC_2</type>
<position>100,148</position>
<input>
<ID>N_in0</ID>344 </input>
<input>
<ID>N_in1</ID>189 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>238</ID>
<type>HA_JUNC_2</type>
<position>102,148</position>
<input>
<ID>N_in0</ID>343 </input>
<input>
<ID>N_in1</ID>178 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>239</ID>
<type>HA_JUNC_2</type>
<position>102,180.5</position>
<input>
<ID>N_in0</ID>178 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>240</ID>
<type>HA_JUNC_2</type>
<position>101,148</position>
<input>
<ID>N_in0</ID>342 </input>
<input>
<ID>N_in1</ID>176 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>241</ID>
<type>HA_JUNC_2</type>
<position>101,180.5</position>
<input>
<ID>N_in0</ID>190 </input>
<input>
<ID>N_in1</ID>574 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>242</ID>
<type>HA_JUNC_2</type>
<position>97.5,177.5</position>
<input>
<ID>N_in0</ID>193 </input>
<input>
<ID>N_in1</ID>179 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>243</ID>
<type>HA_JUNC_2</type>
<position>97.5,178.5</position>
<input>
<ID>N_in0</ID>192 </input>
<input>
<ID>N_in1</ID>180 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>244</ID>
<type>BA_NAND2</type>
<position>114,161</position>
<input>
<ID>IN_0</ID>188 </input>
<input>
<ID>IN_1</ID>187 </input>
<output>
<ID>OUT</ID>183 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>245</ID>
<type>BA_NAND2</type>
<position>114,156.5</position>
<input>
<ID>IN_0</ID>176 </input>
<input>
<ID>IN_1</ID>187 </input>
<output>
<ID>OUT</ID>184 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>246</ID>
<type>HA_JUNC_2</type>
<position>124,177.5</position>
<input>
<ID>N_in0</ID>179 </input>
<input>
<ID>N_in1</ID>210 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>247</ID>
<type>HA_JUNC_2</type>
<position>124,178.5</position>
<input>
<ID>N_in0</ID>180 </input>
<input>
<ID>N_in1</ID>209 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>248</ID>
<type>BA_NAND2</type>
<position>114,152</position>
<input>
<ID>IN_0</ID>188 </input>
<input>
<ID>IN_1</ID>176 </input>
<output>
<ID>OUT</ID>185 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>249</ID>
<type>DA_FROM</type>
<position>109.5,166</position>
<input>
<ID>IN_0</ID>181 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>250</ID>
<type>BI_NANDX3</type>
<position>106.5,156.5</position>
<input>
<ID>IN_0</ID>185 </input>
<input>
<ID>IN_1</ID>184 </input>
<input>
<ID>IN_2</ID>183 </input>
<output>
<ID>OUT</ID>186 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>251</ID>
<type>DA_FROM</type>
<position>109.5,164</position>
<input>
<ID>IN_0</ID>182 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Reset</lparam></gate>
<gate>
<ID>252</ID>
<type>HA_JUNC_2</type>
<position>97.5,156.5</position>
<input>
<ID>N_in0</ID>191 </input>
<input>
<ID>N_in1</ID>186 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>253</ID>
<type>AE_SMALL_INVERTER</type>
<position>122.5,154</position>
<input>
<ID>IN_0</ID>178 </input>
<output>
<ID>OUT_0</ID>188 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>254</ID>
<type>HA_JUNC_2</type>
<position>152.5,156.5</position>
<input>
<ID>N_in0</ID>205 </input>
<input>
<ID>N_in1</ID>227 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>255</ID>
<type>AE_DFF_LOW</type>
<position>144.5,169</position>
<input>
<ID>IN_0</ID>195 </input>
<output>
<ID>OUT_0</ID>194 </output>
<input>
<ID>clear</ID>200 </input>
<input>
<ID>clock</ID>199 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>256</ID>
<type>DE_TO</type>
<position>144,175.5</position>
<input>
<ID>IN_0</ID>194 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 0.2</lparam></gate>
<gate>
<ID>257</ID>
<type>AE_MUX_4x1</type>
<position>136.5,171</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>196 </input>
<input>
<ID>IN_2</ID>208 </input>
<input>
<ID>IN_3</ID>207 </input>
<output>
<ID>OUT</ID>195 </output>
<input>
<ID>SEL_0</ID>198 </input>
<input>
<ID>SEL_1</ID>197 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>258</ID>
<type>HA_JUNC_2</type>
<position>128.5,180.5</position>
<input>
<ID>N_in0</ID>194 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>259</ID>
<type>HA_JUNC_2</type>
<position>128.5,148</position>
<input>
<ID>N_in0</ID>354 </input>
<input>
<ID>N_in1</ID>207 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>260</ID>
<type>HA_JUNC_2</type>
<position>130.5,148</position>
<input>
<ID>N_in0</ID>341 </input>
<input>
<ID>N_in1</ID>196 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>261</ID>
<type>HA_JUNC_2</type>
<position>130.5,180.5</position>
<input>
<ID>N_in0</ID>196 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>262</ID>
<type>HA_JUNC_2</type>
<position>129.5,148</position>
<input>
<ID>N_in0</ID>340 </input>
<input>
<ID>N_in1</ID>194 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>263</ID>
<type>HA_JUNC_2</type>
<position>129.5,180.5</position>
<input>
<ID>N_in0</ID>208 </input>
<input>
<ID>N_in1</ID>574 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>264</ID>
<type>HA_JUNC_2</type>
<position>126,177.5</position>
<input>
<ID>N_in0</ID>210 </input>
<input>
<ID>N_in1</ID>197 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>265</ID>
<type>HA_JUNC_2</type>
<position>126,178.5</position>
<input>
<ID>N_in0</ID>209 </input>
<input>
<ID>N_in1</ID>198 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>266</ID>
<type>BA_NAND2</type>
<position>142.5,161</position>
<input>
<ID>IN_0</ID>206 </input>
<input>
<ID>IN_1</ID>205 </input>
<output>
<ID>OUT</ID>201 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>267</ID>
<type>BA_NAND2</type>
<position>142.5,156.5</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>205 </input>
<output>
<ID>OUT</ID>202 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>268</ID>
<type>HA_JUNC_2</type>
<position>152.5,177.5</position>
<input>
<ID>N_in0</ID>197 </input>
<input>
<ID>N_in1</ID>229 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>269</ID>
<type>HA_JUNC_2</type>
<position>152.5,178.5</position>
<input>
<ID>N_in0</ID>198 </input>
<input>
<ID>N_in1</ID>228 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>270</ID>
<type>BA_NAND2</type>
<position>142.5,152</position>
<input>
<ID>IN_0</ID>206 </input>
<input>
<ID>IN_1</ID>194 </input>
<output>
<ID>OUT</ID>203 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>271</ID>
<type>DA_FROM</type>
<position>138,166</position>
<input>
<ID>IN_0</ID>199 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>272</ID>
<type>BI_NANDX3</type>
<position>135,156.5</position>
<input>
<ID>IN_0</ID>203 </input>
<input>
<ID>IN_1</ID>202 </input>
<input>
<ID>IN_2</ID>201 </input>
<output>
<ID>OUT</ID>204 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>273</ID>
<type>DA_FROM</type>
<position>138,164</position>
<input>
<ID>IN_0</ID>200 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Reset</lparam></gate>
<gate>
<ID>274</ID>
<type>HA_JUNC_2</type>
<position>126,156.5</position>
<input>
<ID>N_in0</ID>211 </input>
<input>
<ID>N_in1</ID>204 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>275</ID>
<type>AE_SMALL_INVERTER</type>
<position>151,154</position>
<input>
<ID>IN_0</ID>196 </input>
<output>
<ID>OUT_0</ID>206 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>276</ID>
<type>HA_JUNC_2</type>
<position>181,156.5</position>
<input>
<ID>N_in0</ID>223 </input>
<input>
<ID>N_in1</ID>245 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>277</ID>
<type>AE_DFF_LOW</type>
<position>173,169</position>
<input>
<ID>IN_0</ID>213 </input>
<output>
<ID>OUT_0</ID>212 </output>
<input>
<ID>clear</ID>218 </input>
<input>
<ID>clock</ID>217 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>278</ID>
<type>DE_TO</type>
<position>172.5,175.5</position>
<input>
<ID>IN_0</ID>212 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 0.1</lparam></gate>
<gate>
<ID>279</ID>
<type>AE_MUX_4x1</type>
<position>165,171</position>
<input>
<ID>IN_0</ID>212 </input>
<input>
<ID>IN_1</ID>214 </input>
<input>
<ID>IN_2</ID>226 </input>
<input>
<ID>IN_3</ID>225 </input>
<output>
<ID>OUT</ID>213 </output>
<input>
<ID>SEL_0</ID>216 </input>
<input>
<ID>SEL_1</ID>215 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>280</ID>
<type>AA_LABEL</type>
<position>75,187.5</position>
<gparam>LABEL_TEXT Full Sorter Circuit</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>281</ID>
<type>HA_JUNC_2</type>
<position>157,180.5</position>
<input>
<ID>N_in0</ID>212 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>282</ID>
<type>HA_JUNC_2</type>
<position>157,148</position>
<input>
<ID>N_in0</ID>353 </input>
<input>
<ID>N_in1</ID>225 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>283</ID>
<type>HA_JUNC_2</type>
<position>159,148</position>
<input>
<ID>N_in0</ID>352 </input>
<input>
<ID>N_in1</ID>214 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>284</ID>
<type>HA_JUNC_2</type>
<position>159,180.5</position>
<input>
<ID>N_in0</ID>214 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>285</ID>
<type>HA_JUNC_2</type>
<position>158,148</position>
<input>
<ID>N_in0</ID>351 </input>
<input>
<ID>N_in1</ID>212 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>286</ID>
<type>HA_JUNC_2</type>
<position>158,180.5</position>
<input>
<ID>N_in0</ID>226 </input>
<input>
<ID>N_in1</ID>574 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>287</ID>
<type>HA_JUNC_2</type>
<position>154.5,177.5</position>
<input>
<ID>N_in0</ID>229 </input>
<input>
<ID>N_in1</ID>215 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>288</ID>
<type>HA_JUNC_2</type>
<position>154.5,178.5</position>
<input>
<ID>N_in0</ID>228 </input>
<input>
<ID>N_in1</ID>216 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>289</ID>
<type>BA_NAND2</type>
<position>171,161</position>
<input>
<ID>IN_0</ID>224 </input>
<input>
<ID>IN_1</ID>223 </input>
<output>
<ID>OUT</ID>219 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>290</ID>
<type>BA_NAND2</type>
<position>171,156.5</position>
<input>
<ID>IN_0</ID>212 </input>
<input>
<ID>IN_1</ID>223 </input>
<output>
<ID>OUT</ID>220 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>291</ID>
<type>HA_JUNC_2</type>
<position>181,177.5</position>
<input>
<ID>N_in0</ID>215 </input>
<input>
<ID>N_in1</ID>247 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>292</ID>
<type>HA_JUNC_2</type>
<position>181,178.5</position>
<input>
<ID>N_in0</ID>216 </input>
<input>
<ID>N_in1</ID>246 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>293</ID>
<type>BA_NAND2</type>
<position>171,152</position>
<input>
<ID>IN_0</ID>224 </input>
<input>
<ID>IN_1</ID>212 </input>
<output>
<ID>OUT</ID>221 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>294</ID>
<type>DA_FROM</type>
<position>166.5,166</position>
<input>
<ID>IN_0</ID>217 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>295</ID>
<type>HA_JUNC_2</type>
<position>81,180.5</position>
<input>
<ID>N_in0</ID>256 </input>
<input>
<ID>N_in1</ID>571 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>296</ID>
<type>BI_NANDX3</type>
<position>163.5,156.5</position>
<input>
<ID>IN_0</ID>221 </input>
<input>
<ID>IN_1</ID>220 </input>
<input>
<ID>IN_2</ID>219 </input>
<output>
<ID>OUT</ID>222 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>297</ID>
<type>HA_JUNC_2</type>
<position>81,148</position>
<input>
<ID>N_in0</ID>350 </input>
<input>
<ID>N_in1</ID>252 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>298</ID>
<type>DA_FROM</type>
<position>166.5,164</position>
<input>
<ID>IN_0</ID>218 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Reset</lparam></gate>
<gate>
<ID>299</ID>
<type>HA_JUNC_2</type>
<position>95.5,178.5</position>
<input>
<ID>N_in0</ID>254 </input>
<input>
<ID>N_in1</ID>192 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>300</ID>
<type>HA_JUNC_2</type>
<position>154.5,156.5</position>
<input>
<ID>N_in0</ID>227 </input>
<input>
<ID>N_in1</ID>222 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>301</ID>
<type>HA_JUNC_2</type>
<position>95.5,177.5</position>
<input>
<ID>N_in0</ID>255 </input>
<input>
<ID>N_in1</ID>193 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>302</ID>
<type>AE_SMALL_INVERTER</type>
<position>179.5,154</position>
<input>
<ID>IN_0</ID>214 </input>
<output>
<ID>OUT_0</ID>224 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>303</ID>
<type>HA_JUNC_2</type>
<position>95.5,156.5</position>
<input>
<ID>N_in0</ID>252 </input>
<input>
<ID>N_in1</ID>191 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>304</ID>
<type>HA_JUNC_2</type>
<position>209.5,156.5</position>
<input>
<ID>N_in0</ID>241 </input>
<input>
<ID>N_in1</ID>248 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>305</ID>
<type>HA_JUNC_2</type>
<position>80,180.5</position>
<input>
<ID>N_in0</ID>251 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>306</ID>
<type>AE_DFF_LOW</type>
<position>201.5,169</position>
<input>
<ID>IN_0</ID>231 </input>
<output>
<ID>OUT_0</ID>230 </output>
<input>
<ID>clear</ID>236 </input>
<input>
<ID>clock</ID>235 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>307</ID>
<type>HA_JUNC_2</type>
<position>80,148</position>
<input>
<ID>N_in0</ID>349 </input>
<input>
<ID>N_in1</ID>251 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>308</ID>
<type>DE_TO</type>
<position>201,175.5</position>
<input>
<ID>IN_0</ID>230 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 0.0</lparam></gate>
<gate>
<ID>309</ID>
<type>AE_MUX_4x1</type>
<position>193.5,171</position>
<input>
<ID>IN_0</ID>230 </input>
<input>
<ID>IN_1</ID>232 </input>
<input>
<ID>IN_2</ID>244 </input>
<input>
<ID>IN_3</ID>243 </input>
<output>
<ID>OUT</ID>231 </output>
<input>
<ID>SEL_0</ID>234 </input>
<input>
<ID>SEL_1</ID>233 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>310</ID>
<type>HA_JUNC_2</type>
<position>185.5,180.5</position>
<input>
<ID>N_in0</ID>230 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>311</ID>
<type>HA_JUNC_2</type>
<position>185.5,148</position>
<input>
<ID>N_in0</ID>348 </input>
<input>
<ID>N_in1</ID>243 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>312</ID>
<type>HA_JUNC_2</type>
<position>187.5,148</position>
<input>
<ID>N_in0</ID>347 </input>
<input>
<ID>N_in1</ID>232 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>313</ID>
<type>AO_XNOR2</type>
<position>84.5,175.5</position>
<input>
<ID>IN_0</ID>256 </input>
<input>
<ID>IN_1</ID>252 </input>
<output>
<ID>OUT</ID>253 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>314</ID>
<type>HA_JUNC_2</type>
<position>187.5,180.5</position>
<input>
<ID>N_in0</ID>232 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>315</ID>
<type>BI_NANDX2</type>
<position>90.5,173</position>
<input>
<ID>IN_0</ID>253 </input>
<input>
<ID>IN_1</ID>257 </input>
<output>
<ID>OUT</ID>254 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>316</ID>
<type>HA_JUNC_2</type>
<position>186.5,113.5</position>
<input>
<ID>N_in0</ID>443 </input>
<input>
<ID>N_in1</ID>312 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>317</ID>
<type>BI_NANDX2</type>
<position>90.5,133.5</position>
<input>
<ID>IN_0</ID>339 </input>
<input>
<ID>IN_1</ID>338 </input>
<output>
<ID>OUT</ID>337 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>318</ID>
<type>HA_JUNC_2</type>
<position>186.5,146</position>
<input>
<ID>N_in0</ID>326 </input>
<input>
<ID>N_in1</ID>346 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>319</ID>
<type>AE_SMALL_INVERTER</type>
<position>83.5,137.5</position>
<input>
<ID>IN_0</ID>333 </input>
<output>
<ID>OUT_0</ID>339 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>320</ID>
<type>HA_JUNC_2</type>
<position>183,143</position>
<input>
<ID>N_in0</ID>329 </input>
<input>
<ID>N_in1</ID>315 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>321</ID>
<type>HA_JUNC_2</type>
<position>183,144</position>
<input>
<ID>N_in0</ID>328 </input>
<input>
<ID>N_in1</ID>316 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>322</ID>
<type>BA_NAND2</type>
<position>199.5,126.5</position>
<input>
<ID>IN_0</ID>324 </input>
<input>
<ID>IN_1</ID>323 </input>
<output>
<ID>OUT</ID>319 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>323</ID>
<type>BA_NAND2</type>
<position>199.5,122</position>
<input>
<ID>IN_0</ID>312 </input>
<input>
<ID>IN_1</ID>323 </input>
<output>
<ID>OUT</ID>320 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>324</ID>
<type>HA_JUNC_2</type>
<position>209.5,143</position>
<input>
<ID>N_in0</ID>315 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>325</ID>
<type>HA_JUNC_2</type>
<position>209.5,144</position>
<input>
<ID>N_in0</ID>316 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>326</ID>
<type>BA_NAND2</type>
<position>199.5,117.5</position>
<input>
<ID>IN_0</ID>324 </input>
<input>
<ID>IN_1</ID>312 </input>
<output>
<ID>OUT</ID>321 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>327</ID>
<type>DA_FROM</type>
<position>195,131.5</position>
<input>
<ID>IN_0</ID>317 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>328</ID>
<type>BI_NANDX3</type>
<position>192,122</position>
<input>
<ID>IN_0</ID>321 </input>
<input>
<ID>IN_1</ID>320 </input>
<input>
<ID>IN_2</ID>319 </input>
<output>
<ID>OUT</ID>322 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>329</ID>
<type>DA_FROM</type>
<position>195,129.5</position>
<input>
<ID>IN_0</ID>318 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Reset</lparam></gate>
<gate>
<ID>330</ID>
<type>HA_JUNC_2</type>
<position>183,122</position>
<input>
<ID>N_in0</ID>327 </input>
<input>
<ID>N_in1</ID>322 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>331</ID>
<type>AE_SMALL_INVERTER</type>
<position>208,119.5</position>
<input>
<ID>IN_0</ID>314 </input>
<output>
<ID>OUT_0</ID>324 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>332</ID>
<type>HA_JUNC_2</type>
<position>211.5,146</position>
<input>
<ID>N_in0</ID>331 </input>
<input>
<ID>N_in1</ID>345 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>333</ID>
<type>HE_JUNC_4</type>
<position>211.5,122</position>
<input>
<ID>N_in0</ID>330 </input>
<input>
<ID>N_in2</ID>332 </input>
<input>
<ID>N_in3</ID>331 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>334</ID>
<type>HA_JUNC_2</type>
<position>211.5,113.5</position>
<input>
<ID>N_in0</ID>442 </input>
<input>
<ID>N_in1</ID>332 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>335</ID>
<type>HA_JUNC_2</type>
<position>124,122</position>
<input>
<ID>N_in0</ID>269 </input>
<input>
<ID>N_in1</ID>293 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>336</ID>
<type>AE_DFF_LOW</type>
<position>116,134.5</position>
<input>
<ID>IN_0</ID>259 </input>
<output>
<ID>OUT_0</ID>258 </output>
<input>
<ID>clear</ID>264 </input>
<input>
<ID>clock</ID>263 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>337</ID>
<type>DE_TO</type>
<position>115.5,141</position>
<input>
<ID>IN_0</ID>258 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1.3</lparam></gate>
<gate>
<ID>338</ID>
<type>AE_MUX_4x1</type>
<position>108,136.5</position>
<input>
<ID>IN_0</ID>258 </input>
<input>
<ID>IN_1</ID>260 </input>
<input>
<ID>IN_2</ID>272 </input>
<input>
<ID>IN_3</ID>271 </input>
<output>
<ID>OUT</ID>259 </output>
<input>
<ID>SEL_0</ID>262 </input>
<input>
<ID>SEL_1</ID>261 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>339</ID>
<type>HA_JUNC_2</type>
<position>100,146</position>
<input>
<ID>N_in0</ID>258 </input>
<input>
<ID>N_in1</ID>344 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>340</ID>
<type>HA_JUNC_2</type>
<position>100,113.5</position>
<input>
<ID>N_in0</ID>441 </input>
<input>
<ID>N_in1</ID>271 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>341</ID>
<type>HA_JUNC_2</type>
<position>102,113.5</position>
<input>
<ID>N_in0</ID>440 </input>
<input>
<ID>N_in1</ID>260 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>342</ID>
<type>HA_JUNC_2</type>
<position>102,146</position>
<input>
<ID>N_in0</ID>260 </input>
<input>
<ID>N_in1</ID>343 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>343</ID>
<type>HA_JUNC_2</type>
<position>101,113.5</position>
<input>
<ID>N_in0</ID>439 </input>
<input>
<ID>N_in1</ID>258 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>344</ID>
<type>HA_JUNC_2</type>
<position>101,146</position>
<input>
<ID>N_in0</ID>272 </input>
<input>
<ID>N_in1</ID>342 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>345</ID>
<type>HA_JUNC_2</type>
<position>97.5,143</position>
<input>
<ID>N_in0</ID>275 </input>
<input>
<ID>N_in1</ID>261 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>346</ID>
<type>HA_JUNC_2</type>
<position>97.5,144</position>
<input>
<ID>N_in0</ID>274 </input>
<input>
<ID>N_in1</ID>262 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>347</ID>
<type>BA_NAND2</type>
<position>114,126.5</position>
<input>
<ID>IN_0</ID>270 </input>
<input>
<ID>IN_1</ID>269 </input>
<output>
<ID>OUT</ID>265 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>348</ID>
<type>BA_NAND2</type>
<position>114,122</position>
<input>
<ID>IN_0</ID>258 </input>
<input>
<ID>IN_1</ID>269 </input>
<output>
<ID>OUT</ID>266 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>349</ID>
<type>HA_JUNC_2</type>
<position>124,143</position>
<input>
<ID>N_in0</ID>261 </input>
<input>
<ID>N_in1</ID>292 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>350</ID>
<type>HA_JUNC_2</type>
<position>124,144</position>
<input>
<ID>N_in0</ID>262 </input>
<input>
<ID>N_in1</ID>291 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>351</ID>
<type>BA_NAND2</type>
<position>114,117.5</position>
<input>
<ID>IN_0</ID>270 </input>
<input>
<ID>IN_1</ID>258 </input>
<output>
<ID>OUT</ID>267 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>352</ID>
<type>DA_FROM</type>
<position>109.5,131.5</position>
<input>
<ID>IN_0</ID>263 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>353</ID>
<type>BI_NANDX3</type>
<position>106.5,122</position>
<input>
<ID>IN_0</ID>267 </input>
<input>
<ID>IN_1</ID>266 </input>
<input>
<ID>IN_2</ID>265 </input>
<output>
<ID>OUT</ID>268 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>354</ID>
<type>DA_FROM</type>
<position>109.5,129.5</position>
<input>
<ID>IN_0</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Reset</lparam></gate>
<gate>
<ID>355</ID>
<type>HA_JUNC_2</type>
<position>97.5,122</position>
<input>
<ID>N_in0</ID>273 </input>
<input>
<ID>N_in1</ID>268 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>356</ID>
<type>AE_SMALL_INVERTER</type>
<position>122.5,119.5</position>
<input>
<ID>IN_0</ID>260 </input>
<output>
<ID>OUT_0</ID>270 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>357</ID>
<type>HA_JUNC_2</type>
<position>152.5,122</position>
<input>
<ID>N_in0</ID>287 </input>
<input>
<ID>N_in1</ID>309 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>358</ID>
<type>AE_DFF_LOW</type>
<position>144.5,134.5</position>
<input>
<ID>IN_0</ID>277 </input>
<output>
<ID>OUT_0</ID>276 </output>
<input>
<ID>clear</ID>282 </input>
<input>
<ID>clock</ID>281 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>359</ID>
<type>DE_TO</type>
<position>144,141</position>
<input>
<ID>IN_0</ID>276 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1.2</lparam></gate>
<gate>
<ID>360</ID>
<type>AE_MUX_4x1</type>
<position>136.5,136.5</position>
<input>
<ID>IN_0</ID>276 </input>
<input>
<ID>IN_1</ID>278 </input>
<input>
<ID>IN_2</ID>290 </input>
<input>
<ID>IN_3</ID>289 </input>
<output>
<ID>OUT</ID>277 </output>
<input>
<ID>SEL_0</ID>280 </input>
<input>
<ID>SEL_1</ID>279 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>361</ID>
<type>HA_JUNC_2</type>
<position>128.5,146</position>
<input>
<ID>N_in0</ID>276 </input>
<input>
<ID>N_in1</ID>354 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>362</ID>
<type>HA_JUNC_2</type>
<position>128.5,113.5</position>
<input>
<ID>N_in0</ID>445 </input>
<input>
<ID>N_in1</ID>289 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>363</ID>
<type>HA_JUNC_2</type>
<position>130.5,113.5</position>
<input>
<ID>N_in0</ID>437 </input>
<input>
<ID>N_in1</ID>278 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>364</ID>
<type>HA_JUNC_2</type>
<position>130.5,146</position>
<input>
<ID>N_in0</ID>278 </input>
<input>
<ID>N_in1</ID>341 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>365</ID>
<type>HA_JUNC_2</type>
<position>129.5,113.5</position>
<input>
<ID>N_in0</ID>438 </input>
<input>
<ID>N_in1</ID>276 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>366</ID>
<type>HA_JUNC_2</type>
<position>129.5,146</position>
<input>
<ID>N_in0</ID>290 </input>
<input>
<ID>N_in1</ID>340 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>367</ID>
<type>HA_JUNC_2</type>
<position>126,143</position>
<input>
<ID>N_in0</ID>292 </input>
<input>
<ID>N_in1</ID>279 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>368</ID>
<type>HA_JUNC_2</type>
<position>126,144</position>
<input>
<ID>N_in0</ID>291 </input>
<input>
<ID>N_in1</ID>280 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>369</ID>
<type>BA_NAND2</type>
<position>142.5,126.5</position>
<input>
<ID>IN_0</ID>288 </input>
<input>
<ID>IN_1</ID>287 </input>
<output>
<ID>OUT</ID>283 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>370</ID>
<type>BA_NAND2</type>
<position>142.5,122</position>
<input>
<ID>IN_0</ID>276 </input>
<input>
<ID>IN_1</ID>287 </input>
<output>
<ID>OUT</ID>284 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>371</ID>
<type>HA_JUNC_2</type>
<position>152.5,143</position>
<input>
<ID>N_in0</ID>279 </input>
<input>
<ID>N_in1</ID>311 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>372</ID>
<type>HA_JUNC_2</type>
<position>152.5,144</position>
<input>
<ID>N_in0</ID>280 </input>
<input>
<ID>N_in1</ID>310 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>373</ID>
<type>BA_NAND2</type>
<position>142.5,117.5</position>
<input>
<ID>IN_0</ID>288 </input>
<input>
<ID>IN_1</ID>276 </input>
<output>
<ID>OUT</ID>285 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>374</ID>
<type>DA_FROM</type>
<position>138,131.5</position>
<input>
<ID>IN_0</ID>281 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>375</ID>
<type>BI_NANDX3</type>
<position>135,122</position>
<input>
<ID>IN_0</ID>285 </input>
<input>
<ID>IN_1</ID>284 </input>
<input>
<ID>IN_2</ID>283 </input>
<output>
<ID>OUT</ID>286 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>376</ID>
<type>DA_FROM</type>
<position>138,129.5</position>
<input>
<ID>IN_0</ID>282 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Reset</lparam></gate>
<gate>
<ID>377</ID>
<type>HA_JUNC_2</type>
<position>126,122</position>
<input>
<ID>N_in0</ID>293 </input>
<input>
<ID>N_in1</ID>286 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>378</ID>
<type>AE_SMALL_INVERTER</type>
<position>151,119.5</position>
<input>
<ID>IN_0</ID>278 </input>
<output>
<ID>OUT_0</ID>288 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>379</ID>
<type>HA_JUNC_2</type>
<position>181,122</position>
<input>
<ID>N_in0</ID>305 </input>
<input>
<ID>N_in1</ID>327 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>380</ID>
<type>AE_DFF_LOW</type>
<position>173,134.5</position>
<input>
<ID>IN_0</ID>295 </input>
<output>
<ID>OUT_0</ID>294 </output>
<input>
<ID>clear</ID>300 </input>
<input>
<ID>clock</ID>299 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>381</ID>
<type>DE_TO</type>
<position>172.5,141</position>
<input>
<ID>IN_0</ID>294 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1.1</lparam></gate>
<gate>
<ID>382</ID>
<type>AE_MUX_4x1</type>
<position>165,136.5</position>
<input>
<ID>IN_0</ID>294 </input>
<input>
<ID>IN_1</ID>296 </input>
<input>
<ID>IN_2</ID>308 </input>
<input>
<ID>IN_3</ID>307 </input>
<output>
<ID>OUT</ID>295 </output>
<input>
<ID>SEL_0</ID>298 </input>
<input>
<ID>SEL_1</ID>297 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>383</ID>
<type>HA_JUNC_2</type>
<position>157,146</position>
<input>
<ID>N_in0</ID>294 </input>
<input>
<ID>N_in1</ID>353 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>384</ID>
<type>HA_JUNC_2</type>
<position>157,113.5</position>
<input>
<ID>N_in0</ID>446 </input>
<input>
<ID>N_in1</ID>307 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>385</ID>
<type>HA_JUNC_2</type>
<position>159,113.5</position>
<input>
<ID>N_in0</ID>447 </input>
<input>
<ID>N_in1</ID>296 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>386</ID>
<type>HA_JUNC_2</type>
<position>159,146</position>
<input>
<ID>N_in0</ID>296 </input>
<input>
<ID>N_in1</ID>352 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>387</ID>
<type>HA_JUNC_2</type>
<position>158,113.5</position>
<input>
<ID>N_in0</ID>444 </input>
<input>
<ID>N_in1</ID>294 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>388</ID>
<type>HA_JUNC_2</type>
<position>158,146</position>
<input>
<ID>N_in0</ID>308 </input>
<input>
<ID>N_in1</ID>351 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>389</ID>
<type>HA_JUNC_2</type>
<position>154.5,143</position>
<input>
<ID>N_in0</ID>311 </input>
<input>
<ID>N_in1</ID>297 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>390</ID>
<type>HA_JUNC_2</type>
<position>154.5,144</position>
<input>
<ID>N_in0</ID>310 </input>
<input>
<ID>N_in1</ID>298 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>391</ID>
<type>BA_NAND2</type>
<position>171,126.5</position>
<input>
<ID>IN_0</ID>306 </input>
<input>
<ID>IN_1</ID>305 </input>
<output>
<ID>OUT</ID>301 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>392</ID>
<type>BA_NAND2</type>
<position>171,122</position>
<input>
<ID>IN_0</ID>294 </input>
<input>
<ID>IN_1</ID>305 </input>
<output>
<ID>OUT</ID>302 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>393</ID>
<type>HA_JUNC_2</type>
<position>181,143</position>
<input>
<ID>N_in0</ID>297 </input>
<input>
<ID>N_in1</ID>329 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>394</ID>
<type>HA_JUNC_2</type>
<position>181,144</position>
<input>
<ID>N_in0</ID>298 </input>
<input>
<ID>N_in1</ID>328 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>395</ID>
<type>BA_NAND2</type>
<position>171,117.5</position>
<input>
<ID>IN_0</ID>306 </input>
<input>
<ID>IN_1</ID>294 </input>
<output>
<ID>OUT</ID>303 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>396</ID>
<type>DA_FROM</type>
<position>166.5,131.5</position>
<input>
<ID>IN_0</ID>299 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>397</ID>
<type>HA_JUNC_2</type>
<position>81,146</position>
<input>
<ID>N_in0</ID>338 </input>
<input>
<ID>N_in1</ID>350 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>398</ID>
<type>BI_NANDX3</type>
<position>163.5,122</position>
<input>
<ID>IN_0</ID>303 </input>
<input>
<ID>IN_1</ID>302 </input>
<input>
<ID>IN_2</ID>301 </input>
<output>
<ID>OUT</ID>304 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>399</ID>
<type>HA_JUNC_2</type>
<position>81,113.5</position>
<input>
<ID>N_in0</ID>450 </input>
<input>
<ID>N_in1</ID>334 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>400</ID>
<type>DA_FROM</type>
<position>166.5,129.5</position>
<input>
<ID>IN_0</ID>300 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Reset</lparam></gate>
<gate>
<ID>401</ID>
<type>HA_JUNC_2</type>
<position>95.5,144</position>
<input>
<ID>N_in0</ID>336 </input>
<input>
<ID>N_in1</ID>274 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>402</ID>
<type>HA_JUNC_2</type>
<position>154.5,122</position>
<input>
<ID>N_in0</ID>309 </input>
<input>
<ID>N_in1</ID>304 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>403</ID>
<type>HA_JUNC_2</type>
<position>95.5,143</position>
<input>
<ID>N_in0</ID>337 </input>
<input>
<ID>N_in1</ID>275 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>404</ID>
<type>AE_SMALL_INVERTER</type>
<position>179.5,119.5</position>
<input>
<ID>IN_0</ID>296 </input>
<output>
<ID>OUT_0</ID>306 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>405</ID>
<type>HA_JUNC_2</type>
<position>95.5,122</position>
<input>
<ID>N_in0</ID>334 </input>
<input>
<ID>N_in1</ID>273 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>406</ID>
<type>HA_JUNC_2</type>
<position>209.5,122</position>
<input>
<ID>N_in0</ID>323 </input>
<input>
<ID>N_in1</ID>330 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>407</ID>
<type>HA_JUNC_2</type>
<position>80,146</position>
<input>
<ID>N_in0</ID>333 </input>
<input>
<ID>N_in1</ID>349 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>408</ID>
<type>AE_DFF_LOW</type>
<position>201.5,134.5</position>
<input>
<ID>IN_0</ID>313 </input>
<output>
<ID>OUT_0</ID>312 </output>
<input>
<ID>clear</ID>318 </input>
<input>
<ID>clock</ID>317 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>409</ID>
<type>HA_JUNC_2</type>
<position>80,113.5</position>
<input>
<ID>N_in0</ID>451 </input>
<input>
<ID>N_in1</ID>333 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>410</ID>
<type>DE_TO</type>
<position>201,141</position>
<input>
<ID>IN_0</ID>312 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1.0</lparam></gate>
<gate>
<ID>411</ID>
<type>AE_MUX_4x1</type>
<position>193.5,136.5</position>
<input>
<ID>IN_0</ID>312 </input>
<input>
<ID>IN_1</ID>314 </input>
<input>
<ID>IN_2</ID>326 </input>
<input>
<ID>IN_3</ID>325 </input>
<output>
<ID>OUT</ID>313 </output>
<input>
<ID>SEL_0</ID>316 </input>
<input>
<ID>SEL_1</ID>315 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>412</ID>
<type>HA_JUNC_2</type>
<position>185.5,146</position>
<input>
<ID>N_in0</ID>312 </input>
<input>
<ID>N_in1</ID>348 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>413</ID>
<type>HA_JUNC_2</type>
<position>185.5,113.5</position>
<input>
<ID>N_in0</ID>448 </input>
<input>
<ID>N_in1</ID>325 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>414</ID>
<type>HA_JUNC_2</type>
<position>187.5,113.5</position>
<input>
<ID>N_in0</ID>449 </input>
<input>
<ID>N_in1</ID>314 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>415</ID>
<type>AO_XNOR2</type>
<position>84.5,141</position>
<input>
<ID>IN_0</ID>338 </input>
<input>
<ID>IN_1</ID>334 </input>
<output>
<ID>OUT</ID>335 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>416</ID>
<type>HA_JUNC_2</type>
<position>187.5,146</position>
<input>
<ID>N_in0</ID>314 </input>
<input>
<ID>N_in1</ID>347 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>417</ID>
<type>BI_NANDX2</type>
<position>90.5,138.5</position>
<input>
<ID>IN_0</ID>335 </input>
<input>
<ID>IN_1</ID>339 </input>
<output>
<ID>OUT</ID>336 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>418</ID>
<type>HA_JUNC_2</type>
<position>186.5,79</position>
<input>
<ID>N_in0</ID>557 </input>
<input>
<ID>N_in1</ID>409 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>419</ID>
<type>BI_NANDX2</type>
<position>90.5,99</position>
<input>
<ID>IN_0</ID>436 </input>
<input>
<ID>IN_1</ID>435 </input>
<output>
<ID>OUT</ID>434 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>420</ID>
<type>HA_JUNC_2</type>
<position>186.5,111.5</position>
<input>
<ID>N_in0</ID>423 </input>
<input>
<ID>N_in1</ID>443 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>421</ID>
<type>AE_SMALL_INVERTER</type>
<position>83.5,103</position>
<input>
<ID>IN_0</ID>430 </input>
<output>
<ID>OUT_0</ID>436 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>422</ID>
<type>HA_JUNC_2</type>
<position>183,108.5</position>
<input>
<ID>N_in0</ID>426 </input>
<input>
<ID>N_in1</ID>412 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>423</ID>
<type>HA_JUNC_2</type>
<position>183,109.5</position>
<input>
<ID>N_in0</ID>425 </input>
<input>
<ID>N_in1</ID>413 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>424</ID>
<type>BA_NAND2</type>
<position>199.5,92</position>
<input>
<ID>IN_0</ID>421 </input>
<input>
<ID>IN_1</ID>420 </input>
<output>
<ID>OUT</ID>416 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>425</ID>
<type>BA_NAND2</type>
<position>199.5,87.5</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>420 </input>
<output>
<ID>OUT</ID>417 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>426</ID>
<type>HA_JUNC_2</type>
<position>209.5,108.5</position>
<input>
<ID>N_in0</ID>412 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>427</ID>
<type>HA_JUNC_2</type>
<position>209.5,109.5</position>
<input>
<ID>N_in0</ID>413 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>428</ID>
<type>BA_NAND2</type>
<position>199.5,83</position>
<input>
<ID>IN_0</ID>421 </input>
<input>
<ID>IN_1</ID>409 </input>
<output>
<ID>OUT</ID>418 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>429</ID>
<type>DA_FROM</type>
<position>195,97</position>
<input>
<ID>IN_0</ID>414 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>430</ID>
<type>BI_NANDX3</type>
<position>192,87.5</position>
<input>
<ID>IN_0</ID>418 </input>
<input>
<ID>IN_1</ID>417 </input>
<input>
<ID>IN_2</ID>416 </input>
<output>
<ID>OUT</ID>419 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>431</ID>
<type>DA_FROM</type>
<position>195,95</position>
<input>
<ID>IN_0</ID>415 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Reset</lparam></gate>
<gate>
<ID>432</ID>
<type>HA_JUNC_2</type>
<position>183,87.5</position>
<input>
<ID>N_in0</ID>424 </input>
<input>
<ID>N_in1</ID>419 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>433</ID>
<type>AE_SMALL_INVERTER</type>
<position>208,85</position>
<input>
<ID>IN_0</ID>411 </input>
<output>
<ID>OUT_0</ID>421 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>434</ID>
<type>HA_JUNC_2</type>
<position>211.5,111.5</position>
<input>
<ID>N_in0</ID>428 </input>
<input>
<ID>N_in1</ID>442 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>435</ID>
<type>HE_JUNC_4</type>
<position>211.5,87.5</position>
<input>
<ID>N_in0</ID>427 </input>
<input>
<ID>N_in2</ID>429 </input>
<input>
<ID>N_in3</ID>428 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>436</ID>
<type>HA_JUNC_2</type>
<position>211.5,79</position>
<input>
<ID>N_in0</ID>556 </input>
<input>
<ID>N_in1</ID>429 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>437</ID>
<type>HA_JUNC_2</type>
<position>124,87.5</position>
<input>
<ID>N_in0</ID>366 </input>
<input>
<ID>N_in1</ID>390 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>438</ID>
<type>AE_DFF_LOW</type>
<position>116,100</position>
<input>
<ID>IN_0</ID>356 </input>
<output>
<ID>OUT_0</ID>355 </output>
<input>
<ID>clear</ID>361 </input>
<input>
<ID>clock</ID>360 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>439</ID>
<type>DE_TO</type>
<position>115.5,106.5</position>
<input>
<ID>IN_0</ID>355 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 2.3</lparam></gate>
<gate>
<ID>440</ID>
<type>AE_MUX_4x1</type>
<position>108,102</position>
<input>
<ID>IN_0</ID>355 </input>
<input>
<ID>IN_1</ID>357 </input>
<input>
<ID>IN_2</ID>369 </input>
<input>
<ID>IN_3</ID>368 </input>
<output>
<ID>OUT</ID>356 </output>
<input>
<ID>SEL_0</ID>359 </input>
<input>
<ID>SEL_1</ID>358 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>441</ID>
<type>HA_JUNC_2</type>
<position>100,111.5</position>
<input>
<ID>N_in0</ID>355 </input>
<input>
<ID>N_in1</ID>441 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>442</ID>
<type>HA_JUNC_2</type>
<position>100,79</position>
<input>
<ID>N_in0</ID>558 </input>
<input>
<ID>N_in1</ID>368 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>443</ID>
<type>HA_JUNC_2</type>
<position>102,79</position>
<input>
<ID>N_in0</ID>560 </input>
<input>
<ID>N_in1</ID>357 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>444</ID>
<type>HA_JUNC_2</type>
<position>102,111.5</position>
<input>
<ID>N_in0</ID>357 </input>
<input>
<ID>N_in1</ID>440 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>445</ID>
<type>HA_JUNC_2</type>
<position>101,79</position>
<input>
<ID>N_in0</ID>561 </input>
<input>
<ID>N_in1</ID>355 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>446</ID>
<type>HA_JUNC_2</type>
<position>101,111.5</position>
<input>
<ID>N_in0</ID>369 </input>
<input>
<ID>N_in1</ID>439 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>447</ID>
<type>HA_JUNC_2</type>
<position>97.5,108.5</position>
<input>
<ID>N_in0</ID>372 </input>
<input>
<ID>N_in1</ID>358 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>448</ID>
<type>HA_JUNC_2</type>
<position>97.5,109.5</position>
<input>
<ID>N_in0</ID>371 </input>
<input>
<ID>N_in1</ID>359 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>449</ID>
<type>BA_NAND2</type>
<position>114,92</position>
<input>
<ID>IN_0</ID>367 </input>
<input>
<ID>IN_1</ID>366 </input>
<output>
<ID>OUT</ID>362 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>450</ID>
<type>BA_NAND2</type>
<position>114,87.5</position>
<input>
<ID>IN_0</ID>355 </input>
<input>
<ID>IN_1</ID>366 </input>
<output>
<ID>OUT</ID>363 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>451</ID>
<type>HA_JUNC_2</type>
<position>124,108.5</position>
<input>
<ID>N_in0</ID>358 </input>
<input>
<ID>N_in1</ID>389 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>452</ID>
<type>HA_JUNC_2</type>
<position>124,109.5</position>
<input>
<ID>N_in0</ID>359 </input>
<input>
<ID>N_in1</ID>388 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>453</ID>
<type>BA_NAND2</type>
<position>114,83</position>
<input>
<ID>IN_0</ID>367 </input>
<input>
<ID>IN_1</ID>355 </input>
<output>
<ID>OUT</ID>364 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>454</ID>
<type>DA_FROM</type>
<position>109.5,97</position>
<input>
<ID>IN_0</ID>360 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>455</ID>
<type>BI_NANDX3</type>
<position>106.5,87.5</position>
<input>
<ID>IN_0</ID>364 </input>
<input>
<ID>IN_1</ID>363 </input>
<input>
<ID>IN_2</ID>362 </input>
<output>
<ID>OUT</ID>365 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>456</ID>
<type>DA_FROM</type>
<position>109.5,95</position>
<input>
<ID>IN_0</ID>361 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Reset</lparam></gate>
<gate>
<ID>457</ID>
<type>HA_JUNC_2</type>
<position>97.5,87.5</position>
<input>
<ID>N_in0</ID>370 </input>
<input>
<ID>N_in1</ID>365 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>458</ID>
<type>AE_SMALL_INVERTER</type>
<position>122.5,85</position>
<input>
<ID>IN_0</ID>357 </input>
<output>
<ID>OUT_0</ID>367 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>459</ID>
<type>HA_JUNC_2</type>
<position>152.5,87.5</position>
<input>
<ID>N_in0</ID>384 </input>
<input>
<ID>N_in1</ID>406 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>460</ID>
<type>AE_DFF_LOW</type>
<position>144.5,100</position>
<input>
<ID>IN_0</ID>374 </input>
<output>
<ID>OUT_0</ID>373 </output>
<input>
<ID>clear</ID>379 </input>
<input>
<ID>clock</ID>378 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>461</ID>
<type>DE_TO</type>
<position>144,106.5</position>
<input>
<ID>IN_0</ID>373 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 2.2</lparam></gate>
<gate>
<ID>462</ID>
<type>AE_MUX_4x1</type>
<position>136.5,102</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>375 </input>
<input>
<ID>IN_2</ID>387 </input>
<input>
<ID>IN_3</ID>386 </input>
<output>
<ID>OUT</ID>374 </output>
<input>
<ID>SEL_0</ID>377 </input>
<input>
<ID>SEL_1</ID>376 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>463</ID>
<type>HA_JUNC_2</type>
<position>128.5,111.5</position>
<input>
<ID>N_in0</ID>373 </input>
<input>
<ID>N_in1</ID>445 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>464</ID>
<type>HA_JUNC_2</type>
<position>128.5,79</position>
<input>
<ID>N_in0</ID>559 </input>
<input>
<ID>N_in1</ID>386 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>465</ID>
<type>HA_JUNC_2</type>
<position>130.5,79</position>
<input>
<ID>N_in0</ID>562 </input>
<input>
<ID>N_in1</ID>375 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>466</ID>
<type>HA_JUNC_2</type>
<position>130.5,111.5</position>
<input>
<ID>N_in0</ID>375 </input>
<input>
<ID>N_in1</ID>437 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>467</ID>
<type>HA_JUNC_2</type>
<position>129.5,79</position>
<input>
<ID>N_in0</ID>563 </input>
<input>
<ID>N_in1</ID>373 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>468</ID>
<type>HA_JUNC_2</type>
<position>129.5,111.5</position>
<input>
<ID>N_in0</ID>387 </input>
<input>
<ID>N_in1</ID>438 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>469</ID>
<type>HA_JUNC_2</type>
<position>126,108.5</position>
<input>
<ID>N_in0</ID>389 </input>
<input>
<ID>N_in1</ID>376 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>470</ID>
<type>HA_JUNC_2</type>
<position>126,109.5</position>
<input>
<ID>N_in0</ID>388 </input>
<input>
<ID>N_in1</ID>377 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>471</ID>
<type>BA_NAND2</type>
<position>142.5,92</position>
<input>
<ID>IN_0</ID>385 </input>
<input>
<ID>IN_1</ID>384 </input>
<output>
<ID>OUT</ID>380 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>472</ID>
<type>BA_NAND2</type>
<position>142.5,87.5</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>384 </input>
<output>
<ID>OUT</ID>381 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>473</ID>
<type>HA_JUNC_2</type>
<position>152.5,108.5</position>
<input>
<ID>N_in0</ID>376 </input>
<input>
<ID>N_in1</ID>408 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>474</ID>
<type>HA_JUNC_2</type>
<position>152.5,109.5</position>
<input>
<ID>N_in0</ID>377 </input>
<input>
<ID>N_in1</ID>407 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>475</ID>
<type>BA_NAND2</type>
<position>142.5,83</position>
<input>
<ID>IN_0</ID>385 </input>
<input>
<ID>IN_1</ID>373 </input>
<output>
<ID>OUT</ID>382 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>476</ID>
<type>DA_FROM</type>
<position>138,97</position>
<input>
<ID>IN_0</ID>378 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>477</ID>
<type>BI_NANDX3</type>
<position>135,87.5</position>
<input>
<ID>IN_0</ID>382 </input>
<input>
<ID>IN_1</ID>381 </input>
<input>
<ID>IN_2</ID>380 </input>
<output>
<ID>OUT</ID>383 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>478</ID>
<type>DA_FROM</type>
<position>138,95</position>
<input>
<ID>IN_0</ID>379 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Reset</lparam></gate>
<gate>
<ID>479</ID>
<type>HA_JUNC_2</type>
<position>126,87.5</position>
<input>
<ID>N_in0</ID>390 </input>
<input>
<ID>N_in1</ID>383 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>480</ID>
<type>AE_SMALL_INVERTER</type>
<position>151,85</position>
<input>
<ID>IN_0</ID>375 </input>
<output>
<ID>OUT_0</ID>385 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>481</ID>
<type>HA_JUNC_2</type>
<position>181,87.5</position>
<input>
<ID>N_in0</ID>402 </input>
<input>
<ID>N_in1</ID>424 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>482</ID>
<type>AE_DFF_LOW</type>
<position>173,100</position>
<input>
<ID>IN_0</ID>392 </input>
<output>
<ID>OUT_0</ID>391 </output>
<input>
<ID>clear</ID>397 </input>
<input>
<ID>clock</ID>396 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>483</ID>
<type>DE_TO</type>
<position>172.5,106.5</position>
<input>
<ID>IN_0</ID>391 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 2.1</lparam></gate>
<gate>
<ID>484</ID>
<type>AE_MUX_4x1</type>
<position>165,102</position>
<input>
<ID>IN_0</ID>391 </input>
<input>
<ID>IN_1</ID>393 </input>
<input>
<ID>IN_2</ID>405 </input>
<input>
<ID>IN_3</ID>404 </input>
<output>
<ID>OUT</ID>392 </output>
<input>
<ID>SEL_0</ID>395 </input>
<input>
<ID>SEL_1</ID>394 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>485</ID>
<type>HA_JUNC_2</type>
<position>157,111.5</position>
<input>
<ID>N_in0</ID>391 </input>
<input>
<ID>N_in1</ID>446 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>486</ID>
<type>HA_JUNC_2</type>
<position>157,79</position>
<input>
<ID>N_in0</ID>564 </input>
<input>
<ID>N_in1</ID>404 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>487</ID>
<type>HA_JUNC_2</type>
<position>159,79</position>
<input>
<ID>N_in0</ID>565 </input>
<input>
<ID>N_in1</ID>393 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>488</ID>
<type>HA_JUNC_2</type>
<position>159,111.5</position>
<input>
<ID>N_in0</ID>393 </input>
<input>
<ID>N_in1</ID>447 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>489</ID>
<type>HA_JUNC_2</type>
<position>158,79</position>
<input>
<ID>N_in0</ID>566 </input>
<input>
<ID>N_in1</ID>391 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>490</ID>
<type>HA_JUNC_2</type>
<position>158,111.5</position>
<input>
<ID>N_in0</ID>405 </input>
<input>
<ID>N_in1</ID>444 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>491</ID>
<type>HA_JUNC_2</type>
<position>154.5,108.5</position>
<input>
<ID>N_in0</ID>408 </input>
<input>
<ID>N_in1</ID>394 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>492</ID>
<type>HA_JUNC_2</type>
<position>154.5,109.5</position>
<input>
<ID>N_in0</ID>407 </input>
<input>
<ID>N_in1</ID>395 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>493</ID>
<type>BA_NAND2</type>
<position>171,92</position>
<input>
<ID>IN_0</ID>403 </input>
<input>
<ID>IN_1</ID>402 </input>
<output>
<ID>OUT</ID>398 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>494</ID>
<type>BA_NAND2</type>
<position>171,87.5</position>
<input>
<ID>IN_0</ID>391 </input>
<input>
<ID>IN_1</ID>402 </input>
<output>
<ID>OUT</ID>399 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>495</ID>
<type>HA_JUNC_2</type>
<position>181,108.5</position>
<input>
<ID>N_in0</ID>394 </input>
<input>
<ID>N_in1</ID>426 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>496</ID>
<type>HA_JUNC_2</type>
<position>181,109.5</position>
<input>
<ID>N_in0</ID>395 </input>
<input>
<ID>N_in1</ID>425 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>497</ID>
<type>BA_NAND2</type>
<position>171,83</position>
<input>
<ID>IN_0</ID>403 </input>
<input>
<ID>IN_1</ID>391 </input>
<output>
<ID>OUT</ID>400 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>498</ID>
<type>DA_FROM</type>
<position>166.5,97</position>
<input>
<ID>IN_0</ID>396 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>499</ID>
<type>HA_JUNC_2</type>
<position>81,111.5</position>
<input>
<ID>N_in0</ID>435 </input>
<input>
<ID>N_in1</ID>450 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>500</ID>
<type>BI_NANDX3</type>
<position>163.5,87.5</position>
<input>
<ID>IN_0</ID>400 </input>
<input>
<ID>IN_1</ID>399 </input>
<input>
<ID>IN_2</ID>398 </input>
<output>
<ID>OUT</ID>401 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>501</ID>
<type>HA_JUNC_2</type>
<position>81,79</position>
<input>
<ID>N_in0</ID>567 </input>
<input>
<ID>N_in1</ID>431 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>502</ID>
<type>DA_FROM</type>
<position>166.5,95</position>
<input>
<ID>IN_0</ID>397 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Reset</lparam></gate>
<gate>
<ID>503</ID>
<type>HA_JUNC_2</type>
<position>95.5,109.5</position>
<input>
<ID>N_in0</ID>433 </input>
<input>
<ID>N_in1</ID>371 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>504</ID>
<type>HA_JUNC_2</type>
<position>154.5,87.5</position>
<input>
<ID>N_in0</ID>406 </input>
<input>
<ID>N_in1</ID>401 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>505</ID>
<type>HA_JUNC_2</type>
<position>95.5,108.5</position>
<input>
<ID>N_in0</ID>434 </input>
<input>
<ID>N_in1</ID>372 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>506</ID>
<type>AE_SMALL_INVERTER</type>
<position>179.5,85</position>
<input>
<ID>IN_0</ID>393 </input>
<output>
<ID>OUT_0</ID>403 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>507</ID>
<type>HA_JUNC_2</type>
<position>95.5,87.5</position>
<input>
<ID>N_in0</ID>431 </input>
<input>
<ID>N_in1</ID>370 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>508</ID>
<type>HA_JUNC_2</type>
<position>209.5,87.5</position>
<input>
<ID>N_in0</ID>420 </input>
<input>
<ID>N_in1</ID>427 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>509</ID>
<type>HA_JUNC_2</type>
<position>80,111.5</position>
<input>
<ID>N_in0</ID>430 </input>
<input>
<ID>N_in1</ID>451 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>510</ID>
<type>AE_DFF_LOW</type>
<position>201.5,100</position>
<input>
<ID>IN_0</ID>410 </input>
<output>
<ID>OUT_0</ID>409 </output>
<input>
<ID>clear</ID>415 </input>
<input>
<ID>clock</ID>414 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>511</ID>
<type>HA_JUNC_2</type>
<position>80,79</position>
<input>
<ID>N_in0</ID>568 </input>
<input>
<ID>N_in1</ID>430 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>512</ID>
<type>DE_TO</type>
<position>201,106.5</position>
<input>
<ID>IN_0</ID>409 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 2.0</lparam></gate>
<gate>
<ID>513</ID>
<type>AE_MUX_4x1</type>
<position>193.5,102</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>411 </input>
<input>
<ID>IN_2</ID>423 </input>
<input>
<ID>IN_3</ID>422 </input>
<output>
<ID>OUT</ID>410 </output>
<input>
<ID>SEL_0</ID>413 </input>
<input>
<ID>SEL_1</ID>412 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>514</ID>
<type>HA_JUNC_2</type>
<position>185.5,111.5</position>
<input>
<ID>N_in0</ID>409 </input>
<input>
<ID>N_in1</ID>448 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>515</ID>
<type>HA_JUNC_2</type>
<position>185.5,79</position>
<input>
<ID>N_in0</ID>569 </input>
<input>
<ID>N_in1</ID>422 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>516</ID>
<type>HA_JUNC_2</type>
<position>187.5,79</position>
<input>
<ID>N_in0</ID>570 </input>
<input>
<ID>N_in1</ID>411 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>517</ID>
<type>AO_XNOR2</type>
<position>84.5,106.5</position>
<input>
<ID>IN_0</ID>435 </input>
<input>
<ID>IN_1</ID>431 </input>
<output>
<ID>OUT</ID>432 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>518</ID>
<type>HA_JUNC_2</type>
<position>187.5,111.5</position>
<input>
<ID>N_in0</ID>411 </input>
<input>
<ID>N_in1</ID>449 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>519</ID>
<type>BI_NANDX2</type>
<position>90.5,104</position>
<input>
<ID>IN_0</ID>432 </input>
<input>
<ID>IN_1</ID>436 </input>
<output>
<ID>OUT</ID>433 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>520</ID>
<type>HA_JUNC_2</type>
<position>186.5,44.5</position>
<input>
<ID>N_in1</ID>528 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>521</ID>
<type>BI_NANDX2</type>
<position>90.5,64.5</position>
<input>
<ID>IN_0</ID>555 </input>
<input>
<ID>IN_1</ID>554 </input>
<output>
<ID>OUT</ID>553 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>522</ID>
<type>HA_JUNC_2</type>
<position>186.5,77</position>
<input>
<ID>N_in0</ID>542 </input>
<input>
<ID>N_in1</ID>557 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>523</ID>
<type>AE_SMALL_INVERTER</type>
<position>83.5,68.5</position>
<input>
<ID>IN_0</ID>549 </input>
<output>
<ID>OUT_0</ID>555 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>524</ID>
<type>HA_JUNC_2</type>
<position>183,74</position>
<input>
<ID>N_in0</ID>545 </input>
<input>
<ID>N_in1</ID>531 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>525</ID>
<type>HA_JUNC_2</type>
<position>183,75</position>
<input>
<ID>N_in0</ID>544 </input>
<input>
<ID>N_in1</ID>532 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>526</ID>
<type>BA_NAND2</type>
<position>199.5,57.5</position>
<input>
<ID>IN_0</ID>540 </input>
<input>
<ID>IN_1</ID>539 </input>
<output>
<ID>OUT</ID>535 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>527</ID>
<type>BA_NAND2</type>
<position>199.5,53</position>
<input>
<ID>IN_0</ID>528 </input>
<input>
<ID>IN_1</ID>539 </input>
<output>
<ID>OUT</ID>536 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>528</ID>
<type>HA_JUNC_2</type>
<position>209.5,74</position>
<input>
<ID>N_in0</ID>531 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>529</ID>
<type>HA_JUNC_2</type>
<position>209.5,75</position>
<input>
<ID>N_in0</ID>532 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>530</ID>
<type>BA_NAND2</type>
<position>199.5,48.5</position>
<input>
<ID>IN_0</ID>540 </input>
<input>
<ID>IN_1</ID>528 </input>
<output>
<ID>OUT</ID>537 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>531</ID>
<type>DA_FROM</type>
<position>195,62.5</position>
<input>
<ID>IN_0</ID>533 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>532</ID>
<type>BI_NANDX3</type>
<position>192,53</position>
<input>
<ID>IN_0</ID>537 </input>
<input>
<ID>IN_1</ID>536 </input>
<input>
<ID>IN_2</ID>535 </input>
<output>
<ID>OUT</ID>538 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>533</ID>
<type>DA_FROM</type>
<position>195,60.5</position>
<input>
<ID>IN_0</ID>534 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Reset</lparam></gate>
<gate>
<ID>534</ID>
<type>HA_JUNC_2</type>
<position>183,53</position>
<input>
<ID>N_in0</ID>543 </input>
<input>
<ID>N_in1</ID>538 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>535</ID>
<type>AE_SMALL_INVERTER</type>
<position>208,50.5</position>
<input>
<ID>IN_0</ID>530 </input>
<output>
<ID>OUT_0</ID>540 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>536</ID>
<type>HA_JUNC_2</type>
<position>211.5,77</position>
<input>
<ID>N_in0</ID>547 </input>
<input>
<ID>N_in1</ID>556 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>537</ID>
<type>HE_JUNC_4</type>
<position>211.5,53</position>
<input>
<ID>N_in0</ID>546 </input>
<input>
<ID>N_in2</ID>548 </input>
<input>
<ID>N_in3</ID>547 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>538</ID>
<type>HA_JUNC_2</type>
<position>211.5,44.5</position>
<input>
<ID>N_in0</ID>573 </input>
<input>
<ID>N_in1</ID>548 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>539</ID>
<type>HA_JUNC_2</type>
<position>124,53</position>
<input>
<ID>N_in0</ID>463 </input>
<input>
<ID>N_in1</ID>509 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>540</ID>
<type>AE_DFF_LOW</type>
<position>116,65.5</position>
<input>
<ID>IN_0</ID>453 </input>
<output>
<ID>OUT_0</ID>452 </output>
<input>
<ID>clear</ID>458 </input>
<input>
<ID>clock</ID>457 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>541</ID>
<type>DE_TO</type>
<position>115.5,72</position>
<input>
<ID>IN_0</ID>452 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 3.3</lparam></gate>
<gate>
<ID>542</ID>
<type>AE_MUX_4x1</type>
<position>108,67.5</position>
<input>
<ID>IN_0</ID>452 </input>
<input>
<ID>IN_1</ID>454 </input>
<input>
<ID>IN_2</ID>466 </input>
<input>
<ID>IN_3</ID>465 </input>
<output>
<ID>OUT</ID>453 </output>
<input>
<ID>SEL_0</ID>456 </input>
<input>
<ID>SEL_1</ID>455 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>543</ID>
<type>HA_JUNC_2</type>
<position>100,77</position>
<input>
<ID>N_in0</ID>452 </input>
<input>
<ID>N_in1</ID>558 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>544</ID>
<type>HA_JUNC_2</type>
<position>100,44.5</position>
<input>
<ID>N_in0</ID>573 </input>
<input>
<ID>N_in1</ID>465 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>545</ID>
<type>HA_JUNC_2</type>
<position>102,44.5</position>
<input>
<ID>N_in0</ID>575 </input>
<input>
<ID>N_in1</ID>454 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>546</ID>
<type>HA_JUNC_2</type>
<position>102,77</position>
<input>
<ID>N_in0</ID>454 </input>
<input>
<ID>N_in1</ID>560 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>547</ID>
<type>HA_JUNC_2</type>
<position>101,44.5</position>
<input>
<ID>N_in1</ID>452 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>548</ID>
<type>HA_JUNC_2</type>
<position>101,77</position>
<input>
<ID>N_in0</ID>466 </input>
<input>
<ID>N_in1</ID>561 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>549</ID>
<type>HA_JUNC_2</type>
<position>97.5,74</position>
<input>
<ID>N_in0</ID>469 </input>
<input>
<ID>N_in1</ID>455 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>550</ID>
<type>HA_JUNC_2</type>
<position>97.5,75</position>
<input>
<ID>N_in0</ID>468 </input>
<input>
<ID>N_in1</ID>456 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>551</ID>
<type>BA_NAND2</type>
<position>114,57.5</position>
<input>
<ID>IN_0</ID>464 </input>
<input>
<ID>IN_1</ID>463 </input>
<output>
<ID>OUT</ID>459 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>552</ID>
<type>BA_NAND2</type>
<position>114,53</position>
<input>
<ID>IN_0</ID>452 </input>
<input>
<ID>IN_1</ID>463 </input>
<output>
<ID>OUT</ID>460 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>553</ID>
<type>HA_JUNC_2</type>
<position>124,74</position>
<input>
<ID>N_in0</ID>455 </input>
<input>
<ID>N_in1</ID>508 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>554</ID>
<type>HA_JUNC_2</type>
<position>124,75</position>
<input>
<ID>N_in0</ID>456 </input>
<input>
<ID>N_in1</ID>507 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>555</ID>
<type>BA_NAND2</type>
<position>114,48.5</position>
<input>
<ID>IN_0</ID>464 </input>
<input>
<ID>IN_1</ID>452 </input>
<output>
<ID>OUT</ID>461 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>556</ID>
<type>DA_FROM</type>
<position>109.5,62.5</position>
<input>
<ID>IN_0</ID>457 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>557</ID>
<type>BI_NANDX3</type>
<position>106.5,53</position>
<input>
<ID>IN_0</ID>461 </input>
<input>
<ID>IN_1</ID>460 </input>
<input>
<ID>IN_2</ID>459 </input>
<output>
<ID>OUT</ID>462 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>558</ID>
<type>DA_FROM</type>
<position>109.5,60.5</position>
<input>
<ID>IN_0</ID>458 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Reset</lparam></gate>
<gate>
<ID>559</ID>
<type>HA_JUNC_2</type>
<position>97.5,53</position>
<input>
<ID>N_in0</ID>467 </input>
<input>
<ID>N_in1</ID>462 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>560</ID>
<type>AE_SMALL_INVERTER</type>
<position>122.5,50.5</position>
<input>
<ID>IN_0</ID>454 </input>
<output>
<ID>OUT_0</ID>464 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>561</ID>
<type>HA_JUNC_2</type>
<position>152.5,53</position>
<input>
<ID>N_in0</ID>481 </input>
<input>
<ID>N_in1</ID>525 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>562</ID>
<type>AE_DFF_LOW</type>
<position>144.5,65.5</position>
<input>
<ID>IN_0</ID>471 </input>
<output>
<ID>OUT_0</ID>470 </output>
<input>
<ID>clear</ID>476 </input>
<input>
<ID>clock</ID>475 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>563</ID>
<type>DE_TO</type>
<position>144,72</position>
<input>
<ID>IN_0</ID>470 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 3.2</lparam></gate>
<gate>
<ID>564</ID>
<type>AE_MUX_4x1</type>
<position>136.5,67.5</position>
<input>
<ID>IN_0</ID>470 </input>
<input>
<ID>IN_1</ID>472 </input>
<input>
<ID>IN_2</ID>506 </input>
<input>
<ID>IN_3</ID>483 </input>
<output>
<ID>OUT</ID>471 </output>
<input>
<ID>SEL_0</ID>474 </input>
<input>
<ID>SEL_1</ID>473 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>565</ID>
<type>HA_JUNC_2</type>
<position>128.5,77</position>
<input>
<ID>N_in0</ID>470 </input>
<input>
<ID>N_in1</ID>559 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>566</ID>
<type>HA_JUNC_2</type>
<position>128.5,44.5</position>
<input>
<ID>N_in0</ID>573 </input>
<input>
<ID>N_in1</ID>483 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>567</ID>
<type>HA_JUNC_2</type>
<position>130.5,44.5</position>
<input>
<ID>N_in0</ID>576 </input>
<input>
<ID>N_in1</ID>472 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>568</ID>
<type>HA_JUNC_2</type>
<position>130.5,77</position>
<input>
<ID>N_in0</ID>472 </input>
<input>
<ID>N_in1</ID>562 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>569</ID>
<type>HA_JUNC_2</type>
<position>129.5,44.5</position>
<input>
<ID>N_in1</ID>470 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>570</ID>
<type>HA_JUNC_2</type>
<position>129.5,77</position>
<input>
<ID>N_in0</ID>506 </input>
<input>
<ID>N_in1</ID>563 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>571</ID>
<type>HA_JUNC_2</type>
<position>126,74</position>
<input>
<ID>N_in0</ID>508 </input>
<input>
<ID>N_in1</ID>473 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>572</ID>
<type>HA_JUNC_2</type>
<position>126,75</position>
<input>
<ID>N_in0</ID>507 </input>
<input>
<ID>N_in1</ID>474 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>573</ID>
<type>BA_NAND2</type>
<position>142.5,57.5</position>
<input>
<ID>IN_0</ID>482 </input>
<input>
<ID>IN_1</ID>481 </input>
<output>
<ID>OUT</ID>477 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>574</ID>
<type>BA_NAND2</type>
<position>142.5,53</position>
<input>
<ID>IN_0</ID>470 </input>
<input>
<ID>IN_1</ID>481 </input>
<output>
<ID>OUT</ID>478 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>575</ID>
<type>HA_JUNC_2</type>
<position>152.5,74</position>
<input>
<ID>N_in0</ID>473 </input>
<input>
<ID>N_in1</ID>527 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>576</ID>
<type>HA_JUNC_2</type>
<position>152.5,75</position>
<input>
<ID>N_in0</ID>474 </input>
<input>
<ID>N_in1</ID>526 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>577</ID>
<type>BA_NAND2</type>
<position>142.5,48.5</position>
<input>
<ID>IN_0</ID>482 </input>
<input>
<ID>IN_1</ID>470 </input>
<output>
<ID>OUT</ID>479 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>578</ID>
<type>DA_FROM</type>
<position>138,62.5</position>
<input>
<ID>IN_0</ID>475 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>579</ID>
<type>BI_NANDX3</type>
<position>135,53</position>
<input>
<ID>IN_0</ID>479 </input>
<input>
<ID>IN_1</ID>478 </input>
<input>
<ID>IN_2</ID>477 </input>
<output>
<ID>OUT</ID>480 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>580</ID>
<type>DA_FROM</type>
<position>138,60.5</position>
<input>
<ID>IN_0</ID>476 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Reset</lparam></gate>
<gate>
<ID>581</ID>
<type>HA_JUNC_2</type>
<position>126,53</position>
<input>
<ID>N_in0</ID>509 </input>
<input>
<ID>N_in1</ID>480 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>583</ID>
<type>AE_SMALL_INVERTER</type>
<position>151,50.5</position>
<input>
<ID>IN_0</ID>472 </input>
<output>
<ID>OUT_0</ID>482 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>584</ID>
<type>HA_JUNC_2</type>
<position>181,53</position>
<input>
<ID>N_in0</ID>521 </input>
<input>
<ID>N_in1</ID>543 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>586</ID>
<type>AE_DFF_LOW</type>
<position>173,65.5</position>
<input>
<ID>IN_0</ID>511 </input>
<output>
<ID>OUT_0</ID>510 </output>
<input>
<ID>clear</ID>516 </input>
<input>
<ID>clock</ID>515 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>587</ID>
<type>DE_TO</type>
<position>172.5,72</position>
<input>
<ID>IN_0</ID>510 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 3.1</lparam></gate>
<gate>
<ID>588</ID>
<type>AE_MUX_4x1</type>
<position>165,67.5</position>
<input>
<ID>IN_0</ID>510 </input>
<input>
<ID>IN_1</ID>512 </input>
<input>
<ID>IN_2</ID>524 </input>
<input>
<ID>IN_3</ID>523 </input>
<output>
<ID>OUT</ID>511 </output>
<input>
<ID>SEL_0</ID>514 </input>
<input>
<ID>SEL_1</ID>513 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>589</ID>
<type>HA_JUNC_2</type>
<position>157,77</position>
<input>
<ID>N_in0</ID>510 </input>
<input>
<ID>N_in1</ID>564 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>590</ID>
<type>HA_JUNC_2</type>
<position>157,44.5</position>
<input>
<ID>N_in0</ID>573 </input>
<input>
<ID>N_in1</ID>523 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>591</ID>
<type>HA_JUNC_2</type>
<position>159,44.5</position>
<input>
<ID>N_in0</ID>577 </input>
<input>
<ID>N_in1</ID>512 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>592</ID>
<type>HA_JUNC_2</type>
<position>159,77</position>
<input>
<ID>N_in0</ID>512 </input>
<input>
<ID>N_in1</ID>565 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>593</ID>
<type>HA_JUNC_2</type>
<position>158,44.5</position>
<input>
<ID>N_in1</ID>510 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>594</ID>
<type>HA_JUNC_2</type>
<position>158,77</position>
<input>
<ID>N_in0</ID>524 </input>
<input>
<ID>N_in1</ID>566 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>595</ID>
<type>HA_JUNC_2</type>
<position>154.5,74</position>
<input>
<ID>N_in0</ID>527 </input>
<input>
<ID>N_in1</ID>513 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>596</ID>
<type>HA_JUNC_2</type>
<position>154.5,75</position>
<input>
<ID>N_in0</ID>526 </input>
<input>
<ID>N_in1</ID>514 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>597</ID>
<type>BA_NAND2</type>
<position>171,57.5</position>
<input>
<ID>IN_0</ID>522 </input>
<input>
<ID>IN_1</ID>521 </input>
<output>
<ID>OUT</ID>517 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>598</ID>
<type>BA_NAND2</type>
<position>171,53</position>
<input>
<ID>IN_0</ID>510 </input>
<input>
<ID>IN_1</ID>521 </input>
<output>
<ID>OUT</ID>518 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>599</ID>
<type>HA_JUNC_2</type>
<position>181,74</position>
<input>
<ID>N_in0</ID>513 </input>
<input>
<ID>N_in1</ID>545 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>600</ID>
<type>HA_JUNC_2</type>
<position>181,75</position>
<input>
<ID>N_in0</ID>514 </input>
<input>
<ID>N_in1</ID>544 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>601</ID>
<type>BA_NAND2</type>
<position>171,48.5</position>
<input>
<ID>IN_0</ID>522 </input>
<input>
<ID>IN_1</ID>510 </input>
<output>
<ID>OUT</ID>519 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>602</ID>
<type>DA_FROM</type>
<position>166.5,62.5</position>
<input>
<ID>IN_0</ID>515 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>603</ID>
<type>HA_JUNC_2</type>
<position>81,77</position>
<input>
<ID>N_in0</ID>554 </input>
<input>
<ID>N_in1</ID>567 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>604</ID>
<type>BI_NANDX3</type>
<position>163.5,53</position>
<input>
<ID>IN_0</ID>519 </input>
<input>
<ID>IN_1</ID>518 </input>
<input>
<ID>IN_2</ID>517 </input>
<output>
<ID>OUT</ID>520 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>605</ID>
<type>HA_JUNC_2</type>
<position>81,44.5</position>
<input>
<ID>N_in1</ID>550 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>607</ID>
<type>DA_FROM</type>
<position>166.5,60.5</position>
<input>
<ID>IN_0</ID>516 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Reset</lparam></gate>
<gate>
<ID>608</ID>
<type>HA_JUNC_2</type>
<position>95.5,75</position>
<input>
<ID>N_in0</ID>552 </input>
<input>
<ID>N_in1</ID>468 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>609</ID>
<type>HA_JUNC_2</type>
<position>154.5,53</position>
<input>
<ID>N_in0</ID>525 </input>
<input>
<ID>N_in1</ID>520 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>610</ID>
<type>HA_JUNC_2</type>
<position>95.5,74</position>
<input>
<ID>N_in0</ID>553 </input>
<input>
<ID>N_in1</ID>469 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>612</ID>
<type>AE_SMALL_INVERTER</type>
<position>179.5,50.5</position>
<input>
<ID>IN_0</ID>512 </input>
<output>
<ID>OUT_0</ID>522 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>613</ID>
<type>HA_JUNC_2</type>
<position>95.5,53</position>
<input>
<ID>N_in0</ID>550 </input>
<input>
<ID>N_in1</ID>467 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>614</ID>
<type>HA_JUNC_2</type>
<position>209.5,53</position>
<input>
<ID>N_in0</ID>539 </input>
<input>
<ID>N_in1</ID>546 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>615</ID>
<type>HA_JUNC_2</type>
<position>80,77</position>
<input>
<ID>N_in0</ID>549 </input>
<input>
<ID>N_in1</ID>568 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>616</ID>
<type>AE_DFF_LOW</type>
<position>201.5,65.5</position>
<input>
<ID>IN_0</ID>529 </input>
<output>
<ID>OUT_0</ID>528 </output>
<input>
<ID>clear</ID>534 </input>
<input>
<ID>clock</ID>533 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>617</ID>
<type>HA_JUNC_2</type>
<position>80,44.5</position>
<input>
<ID>N_in0</ID>572 </input>
<input>
<ID>N_in1</ID>549 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>618</ID>
<type>DE_TO</type>
<position>201,72</position>
<input>
<ID>IN_0</ID>528 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 3.0</lparam></gate>
<gate>
<ID>619</ID>
<type>AE_MUX_4x1</type>
<position>193.5,67.5</position>
<input>
<ID>IN_0</ID>528 </input>
<input>
<ID>IN_1</ID>530 </input>
<input>
<ID>IN_2</ID>542 </input>
<input>
<ID>IN_3</ID>541 </input>
<output>
<ID>OUT</ID>529 </output>
<input>
<ID>SEL_0</ID>532 </input>
<input>
<ID>SEL_1</ID>531 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>620</ID>
<type>HA_JUNC_2</type>
<position>185.5,77</position>
<input>
<ID>N_in0</ID>528 </input>
<input>
<ID>N_in1</ID>569 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>621</ID>
<type>HA_JUNC_2</type>
<position>185.5,44.5</position>
<input>
<ID>N_in0</ID>573 </input>
<input>
<ID>N_in1</ID>541 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>622</ID>
<type>HA_JUNC_2</type>
<position>187.5,44.5</position>
<input>
<ID>N_in0</ID>578 </input>
<input>
<ID>N_in1</ID>530 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>624</ID>
<type>AO_XNOR2</type>
<position>84.5,72</position>
<input>
<ID>IN_0</ID>554 </input>
<input>
<ID>IN_1</ID>550 </input>
<output>
<ID>OUT</ID>551 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>625</ID>
<type>HA_JUNC_2</type>
<position>187.5,77</position>
<input>
<ID>N_in0</ID>530 </input>
<input>
<ID>N_in1</ID>570 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>626</ID>
<type>BI_NANDX2</type>
<position>90.5,69.5</position>
<input>
<ID>IN_0</ID>551 </input>
<input>
<ID>IN_1</ID>555 </input>
<output>
<ID>OUT</ID>552 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>628</ID>
<type>EE_VDD</type>
<position>81,183.5</position>
<output>
<ID>OUT_0</ID>571 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>633</ID>
<type>DA_FROM</type>
<position>77,42</position>
<input>
<ID>IN_0</ID>572 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r/w</lparam></gate>
<gate>
<ID>635</ID>
<type>FF_GND</type>
<position>211.5,41.5</position>
<output>
<ID>OUT_0</ID>573 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>636</ID>
<type>DA_FROM</type>
<position>98,39</position>
<input>
<ID>IN_0</ID>575 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>638</ID>
<type>DA_FROM</type>
<position>98,37</position>
<input>
<ID>IN_0</ID>576 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>639</ID>
<type>DA_FROM</type>
<position>98,35</position>
<input>
<ID>IN_0</ID>577 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>640</ID>
<type>DA_FROM</type>
<position>98,33</position>
<input>
<ID>IN_0</ID>578 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<wire>
<ID>389</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,108.5,125,108.5</points>
<connection>
<GID>451</GID>
<name>N_in1</name></connection>
<connection>
<GID>469</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>390</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,87.5,125,87.5</points>
<connection>
<GID>437</GID>
<name>N_in1</name></connection>
<connection>
<GID>479</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177,79.5,177,104.5</points>
<intersection>79.5 2</intersection>
<intersection>84 14</intersection>
<intersection>102 7</intersection>
<intersection>104.5 30</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>157,79.5,177,79.5</points>
<intersection>157 4</intersection>
<intersection>158 17</intersection>
<intersection>177 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>157,79.5,157,110.5</points>
<connection>
<GID>485</GID>
<name>N_in0</name></connection>
<intersection>79.5 2</intersection>
<intersection>99 9</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>176,102,177,102</points>
<connection>
<GID>482</GID>
<name>OUT_0</name></connection>
<intersection>177 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>157,99,162,99</points>
<connection>
<GID>484</GID>
<name>IN_0</name></connection>
<intersection>157 4</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>174,84,177,84</points>
<connection>
<GID>497</GID>
<name>IN_1</name></connection>
<intersection>174 27</intersection>
<intersection>177 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>158,79.5,158,80</points>
<connection>
<GID>489</GID>
<name>N_in1</name></connection>
<intersection>79.5 2</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>174,84,174,86.5</points>
<connection>
<GID>494</GID>
<name>IN_0</name></connection>
<intersection>84 14</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>170.5,104.5,177,104.5</points>
<intersection>170.5 32</intersection>
<intersection>177 0</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>170.5,104.5,170.5,106.5</points>
<connection>
<GID>483</GID>
<name>IN_0</name></connection>
<intersection>104.5 30</intersection></vsegment></shape></wire>
<wire>
<ID>392</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>168,102,170,102</points>
<connection>
<GID>484</GID>
<name>OUT</name></connection>
<connection>
<GID>482</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>393</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,79,159,110.5</points>
<connection>
<GID>488</GID>
<name>N_in0</name></connection>
<connection>
<GID>487</GID>
<name>N_in1</name></connection>
<intersection>79 6</intersection>
<intersection>101 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>159,101,162,101</points>
<connection>
<GID>484</GID>
<name>IN_1</name></connection>
<intersection>159 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>159,79,181.5,79</points>
<intersection>159 0</intersection>
<intersection>181.5 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>181.5,79,181.5,85</points>
<connection>
<GID>506</GID>
<name>IN_0</name></connection>
<intersection>79 6</intersection></vsegment></shape></wire>
<wire>
<ID>394</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165,107,165,108.5</points>
<connection>
<GID>484</GID>
<name>SEL_1</name></connection>
<intersection>108.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>155.5,108.5,180,108.5</points>
<connection>
<GID>495</GID>
<name>N_in0</name></connection>
<connection>
<GID>491</GID>
<name>N_in1</name></connection>
<intersection>165 0</intersection></hsegment></shape></wire>
<wire>
<ID>395</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,107,166,109.5</points>
<connection>
<GID>484</GID>
<name>SEL_0</name></connection>
<intersection>109.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>155.5,109.5,180,109.5</points>
<connection>
<GID>496</GID>
<name>N_in0</name></connection>
<connection>
<GID>492</GID>
<name>N_in1</name></connection>
<intersection>166 0</intersection></hsegment></shape></wire>
<wire>
<ID>396</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,97,170,99</points>
<connection>
<GID>482</GID>
<name>clock</name></connection>
<intersection>97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168.5,97,170,97</points>
<connection>
<GID>498</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment></shape></wire>
<wire>
<ID>397</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173,95,173,96</points>
<connection>
<GID>482</GID>
<name>clear</name></connection>
<intersection>95 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>168.5,95,173,95</points>
<connection>
<GID>502</GID>
<name>IN_0</name></connection>
<intersection>173 0</intersection></hsegment></shape></wire>
<wire>
<ID>398</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,89.5,167,92</points>
<intersection>89.5 1</intersection>
<intersection>92 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166.5,89.5,167,89.5</points>
<connection>
<GID>500</GID>
<name>IN_2</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>167,92,168,92</points>
<connection>
<GID>493</GID>
<name>OUT</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>399</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>166.5,87.5,168,87.5</points>
<connection>
<GID>500</GID>
<name>IN_1</name></connection>
<connection>
<GID>494</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>400</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,83,167,85.5</points>
<intersection>83 1</intersection>
<intersection>85.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167,83,168,83</points>
<connection>
<GID>497</GID>
<name>OUT</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>166.5,85.5,167,85.5</points>
<connection>
<GID>500</GID>
<name>IN_0</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>401</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>155.5,87.5,160.5,87.5</points>
<connection>
<GID>504</GID>
<name>N_in1</name></connection>
<connection>
<GID>500</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>402</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178,87.5,178,93</points>
<intersection>87.5 8</intersection>
<intersection>88.5 1</intersection>
<intersection>93 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>174,88.5,178,88.5</points>
<connection>
<GID>494</GID>
<name>IN_1</name></connection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>174,93,178,93</points>
<connection>
<GID>493</GID>
<name>IN_1</name></connection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>178,87.5,180,87.5</points>
<connection>
<GID>481</GID>
<name>N_in0</name></connection>
<intersection>178 0</intersection></hsegment></shape></wire>
<wire>
<ID>403</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176,82,176,91</points>
<intersection>82 3</intersection>
<intersection>85 2</intersection>
<intersection>91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>174,91,176,91</points>
<connection>
<GID>493</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>176,85,177.5,85</points>
<connection>
<GID>506</GID>
<name>OUT_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>174,82,176,82</points>
<connection>
<GID>497</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment></shape></wire>
<wire>
<ID>404</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,80,156.5,105</points>
<intersection>80 2</intersection>
<intersection>105 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156.5,105,162,105</points>
<connection>
<GID>484</GID>
<name>IN_3</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156.5,80,157,80</points>
<connection>
<GID>486</GID>
<name>N_in1</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>405</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158,103,158,110.5</points>
<connection>
<GID>490</GID>
<name>N_in0</name></connection>
<intersection>103 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>158,103,162,103</points>
<connection>
<GID>484</GID>
<name>IN_2</name></connection>
<intersection>158 0</intersection></hsegment></shape></wire>
<wire>
<ID>406</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153.5,87.5,153.5,87.5</points>
<connection>
<GID>459</GID>
<name>N_in1</name></connection>
<connection>
<GID>504</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>407</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153.5,109.5,153.5,109.5</points>
<connection>
<GID>474</GID>
<name>N_in1</name></connection>
<connection>
<GID>492</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>408</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153.5,108.5,153.5,108.5</points>
<connection>
<GID>473</GID>
<name>N_in1</name></connection>
<connection>
<GID>491</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>409</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205.5,79.5,205.5,104.5</points>
<intersection>79.5 2</intersection>
<intersection>84 14</intersection>
<intersection>102 7</intersection>
<intersection>104.5 30</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>185.5,79.5,205.5,79.5</points>
<intersection>185.5 4</intersection>
<intersection>186.5 17</intersection>
<intersection>205.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>185.5,79.5,185.5,110.5</points>
<connection>
<GID>514</GID>
<name>N_in0</name></connection>
<intersection>79.5 2</intersection>
<intersection>99 9</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>204.5,102,205.5,102</points>
<connection>
<GID>510</GID>
<name>OUT_0</name></connection>
<intersection>205.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>185.5,99,190.5,99</points>
<connection>
<GID>513</GID>
<name>IN_0</name></connection>
<intersection>185.5 4</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>202.5,84,205.5,84</points>
<connection>
<GID>428</GID>
<name>IN_1</name></connection>
<intersection>202.5 27</intersection>
<intersection>205.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>186.5,79.5,186.5,80</points>
<connection>
<GID>418</GID>
<name>N_in1</name></connection>
<intersection>79.5 2</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>202.5,84,202.5,86.5</points>
<connection>
<GID>425</GID>
<name>IN_0</name></connection>
<intersection>84 14</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>199,104.5,205.5,104.5</points>
<intersection>199 32</intersection>
<intersection>205.5 0</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>199,104.5,199,106.5</points>
<connection>
<GID>512</GID>
<name>IN_0</name></connection>
<intersection>104.5 30</intersection></vsegment></shape></wire>
<wire>
<ID>410</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>196.5,102,198.5,102</points>
<connection>
<GID>513</GID>
<name>OUT</name></connection>
<connection>
<GID>510</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>411</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,79,187.5,110.5</points>
<connection>
<GID>518</GID>
<name>N_in0</name></connection>
<connection>
<GID>516</GID>
<name>N_in1</name></connection>
<intersection>79 6</intersection>
<intersection>101 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>187.5,101,190.5,101</points>
<connection>
<GID>513</GID>
<name>IN_1</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>187.5,79,210,79</points>
<intersection>187.5 0</intersection>
<intersection>210 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>210,79,210,85</points>
<connection>
<GID>433</GID>
<name>IN_0</name></connection>
<intersection>79 6</intersection></vsegment></shape></wire>
<wire>
<ID>412</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>193.5,107,193.5,108.5</points>
<connection>
<GID>513</GID>
<name>SEL_1</name></connection>
<intersection>108.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184,108.5,208.5,108.5</points>
<connection>
<GID>426</GID>
<name>N_in0</name></connection>
<connection>
<GID>422</GID>
<name>N_in1</name></connection>
<intersection>193.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>413</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,107,194.5,109.5</points>
<connection>
<GID>513</GID>
<name>SEL_0</name></connection>
<intersection>109.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184,109.5,208.5,109.5</points>
<connection>
<GID>427</GID>
<name>N_in0</name></connection>
<connection>
<GID>423</GID>
<name>N_in1</name></connection>
<intersection>194.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>414</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,97,198.5,99</points>
<connection>
<GID>510</GID>
<name>clock</name></connection>
<intersection>97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>197,97,198.5,97</points>
<connection>
<GID>429</GID>
<name>IN_0</name></connection>
<intersection>198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>415</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201.5,95,201.5,96</points>
<connection>
<GID>510</GID>
<name>clear</name></connection>
<intersection>95 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>197,95,201.5,95</points>
<connection>
<GID>431</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>416</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>195.5,89.5,195.5,92</points>
<intersection>89.5 1</intersection>
<intersection>92 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>195,89.5,195.5,89.5</points>
<connection>
<GID>430</GID>
<name>IN_2</name></connection>
<intersection>195.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>195.5,92,196.5,92</points>
<connection>
<GID>424</GID>
<name>OUT</name></connection>
<intersection>195.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>417</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,87.5,196.5,87.5</points>
<connection>
<GID>430</GID>
<name>IN_1</name></connection>
<connection>
<GID>425</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>418</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>195.5,83,195.5,85.5</points>
<intersection>83 1</intersection>
<intersection>85.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>195.5,83,196.5,83</points>
<connection>
<GID>428</GID>
<name>OUT</name></connection>
<intersection>195.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>195,85.5,195.5,85.5</points>
<connection>
<GID>430</GID>
<name>IN_0</name></connection>
<intersection>195.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>419</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>184,87.5,189,87.5</points>
<connection>
<GID>432</GID>
<name>N_in1</name></connection>
<connection>
<GID>430</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>420</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206.5,87.5,206.5,93</points>
<intersection>87.5 8</intersection>
<intersection>88.5 1</intersection>
<intersection>93 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>202.5,88.5,206.5,88.5</points>
<connection>
<GID>425</GID>
<name>IN_1</name></connection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>202.5,93,206.5,93</points>
<connection>
<GID>424</GID>
<name>IN_1</name></connection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>206.5,87.5,208.5,87.5</points>
<connection>
<GID>508</GID>
<name>N_in0</name></connection>
<intersection>206.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>421</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204.5,82,204.5,91</points>
<intersection>82 3</intersection>
<intersection>85 2</intersection>
<intersection>91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>202.5,91,204.5,91</points>
<connection>
<GID>424</GID>
<name>IN_0</name></connection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>204.5,85,206,85</points>
<connection>
<GID>433</GID>
<name>OUT_0</name></connection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>202.5,82,204.5,82</points>
<connection>
<GID>428</GID>
<name>IN_0</name></connection>
<intersection>204.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>422</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,80,185,105</points>
<intersection>80 2</intersection>
<intersection>105 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185,105,190.5,105</points>
<connection>
<GID>513</GID>
<name>IN_3</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>185,80,185.5,80</points>
<connection>
<GID>515</GID>
<name>N_in1</name></connection>
<intersection>185 0</intersection></hsegment></shape></wire>
<wire>
<ID>423</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186.5,103,186.5,110.5</points>
<connection>
<GID>420</GID>
<name>N_in0</name></connection>
<intersection>103 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>186.5,103,190.5,103</points>
<connection>
<GID>513</GID>
<name>IN_2</name></connection>
<intersection>186.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>424</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182,87.5,182,87.5</points>
<connection>
<GID>432</GID>
<name>N_in0</name></connection>
<connection>
<GID>481</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>425</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182,109.5,182,109.5</points>
<connection>
<GID>423</GID>
<name>N_in0</name></connection>
<connection>
<GID>496</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>426</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182,108.5,182,108.5</points>
<connection>
<GID>422</GID>
<name>N_in0</name></connection>
<connection>
<GID>495</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>427</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210.5,87.5,210.5,87.5</points>
<connection>
<GID>435</GID>
<name>N_in0</name></connection>
<connection>
<GID>508</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>428</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211.5,88.5,211.5,110.5</points>
<connection>
<GID>435</GID>
<name>N_in3</name></connection>
<connection>
<GID>434</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>429</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211.5,80,211.5,86.5</points>
<connection>
<GID>436</GID>
<name>N_in1</name></connection>
<connection>
<GID>435</GID>
<name>N_in2</name></connection></vsegment></shape></wire>
<wire>
<ID>430</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,80,80,110.5</points>
<connection>
<GID>511</GID>
<name>N_in1</name></connection>
<connection>
<GID>509</GID>
<name>N_in0</name></connection>
<intersection>103 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>80,103,81.5,103</points>
<connection>
<GID>421</GID>
<name>IN_0</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>431</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>80.5,87.5,94.5,87.5</points>
<connection>
<GID>507</GID>
<name>N_in0</name></connection>
<intersection>80.5 8</intersection>
<intersection>81 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>81,80,81,87.5</points>
<connection>
<GID>501</GID>
<name>N_in1</name></connection>
<intersection>87.5 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>80.5,87.5,80.5,105.5</points>
<intersection>87.5 2</intersection>
<intersection>105.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>80.5,105.5,81.5,105.5</points>
<connection>
<GID>517</GID>
<name>IN_1</name></connection>
<intersection>80.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>432</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,105,87.5,106.5</points>
<connection>
<GID>519</GID>
<name>IN_0</name></connection>
<connection>
<GID>517</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>433</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,104,93.5,109.5</points>
<connection>
<GID>519</GID>
<name>OUT</name></connection>
<intersection>109.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93.5,109.5,94.5,109.5</points>
<connection>
<GID>503</GID>
<name>N_in0</name></connection>
<intersection>93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>434</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94.5,99,94.5,108.5</points>
<connection>
<GID>505</GID>
<name>N_in0</name></connection>
<intersection>99 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>93.5,99,94.5,99</points>
<connection>
<GID>419</GID>
<name>OUT</name></connection>
<intersection>94.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>435</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,98,81,110.5</points>
<connection>
<GID>499</GID>
<name>N_in0</name></connection>
<intersection>98 3</intersection>
<intersection>107.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81,107.5,81.5,107.5</points>
<connection>
<GID>517</GID>
<name>IN_0</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>81,98,87.5,98</points>
<connection>
<GID>419</GID>
<name>IN_1</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>436</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,103,87.5,103</points>
<connection>
<GID>519</GID>
<name>IN_1</name></connection>
<connection>
<GID>421</GID>
<name>OUT_0</name></connection>
<intersection>86.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>86.5,100,86.5,103</points>
<intersection>100 8</intersection>
<intersection>103 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>86.5,100,87.5,100</points>
<connection>
<GID>419</GID>
<name>IN_0</name></connection>
<intersection>86.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>437</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,112.5,130.5,112.5</points>
<connection>
<GID>363</GID>
<name>N_in0</name></connection>
<connection>
<GID>466</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>438</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,112.5,129.5,112.5</points>
<connection>
<GID>365</GID>
<name>N_in0</name></connection>
<connection>
<GID>468</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>439</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,112.5,101,112.5</points>
<connection>
<GID>343</GID>
<name>N_in0</name></connection>
<connection>
<GID>446</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>440</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,112.5,102,112.5</points>
<connection>
<GID>341</GID>
<name>N_in0</name></connection>
<connection>
<GID>444</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>441</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,112.5,100,112.5</points>
<connection>
<GID>340</GID>
<name>N_in0</name></connection>
<connection>
<GID>441</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>442</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211.5,112.5,211.5,112.5</points>
<connection>
<GID>334</GID>
<name>N_in0</name></connection>
<connection>
<GID>434</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>443</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186.5,112.5,186.5,112.5</points>
<connection>
<GID>316</GID>
<name>N_in0</name></connection>
<connection>
<GID>420</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>444</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158,112.5,158,112.5</points>
<connection>
<GID>387</GID>
<name>N_in0</name></connection>
<connection>
<GID>490</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>445</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128.5,112.5,128.5,112.5</points>
<connection>
<GID>362</GID>
<name>N_in0</name></connection>
<connection>
<GID>463</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>446</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157,112.5,157,112.5</points>
<connection>
<GID>384</GID>
<name>N_in0</name></connection>
<connection>
<GID>485</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>447</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,112.5,159,112.5</points>
<connection>
<GID>385</GID>
<name>N_in0</name></connection>
<connection>
<GID>488</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>448</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185.5,112.5,185.5,112.5</points>
<connection>
<GID>413</GID>
<name>N_in0</name></connection>
<connection>
<GID>514</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>449</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,112.5,187.5,112.5</points>
<connection>
<GID>414</GID>
<name>N_in0</name></connection>
<connection>
<GID>518</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>450</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,112.5,81,112.5</points>
<connection>
<GID>399</GID>
<name>N_in0</name></connection>
<connection>
<GID>499</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>451</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,112.5,80,112.5</points>
<connection>
<GID>409</GID>
<name>N_in0</name></connection>
<connection>
<GID>509</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>452</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,45,120,70</points>
<intersection>45 2</intersection>
<intersection>49.5 14</intersection>
<intersection>67.5 7</intersection>
<intersection>70 30</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>100,45,120,45</points>
<intersection>100 4</intersection>
<intersection>101 17</intersection>
<intersection>120 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>100,45,100,76</points>
<connection>
<GID>543</GID>
<name>N_in0</name></connection>
<intersection>45 2</intersection>
<intersection>64.5 9</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>119,67.5,120,67.5</points>
<connection>
<GID>540</GID>
<name>OUT_0</name></connection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>100,64.5,105,64.5</points>
<connection>
<GID>542</GID>
<name>IN_0</name></connection>
<intersection>100 4</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>117,49.5,120,49.5</points>
<connection>
<GID>555</GID>
<name>IN_1</name></connection>
<intersection>117 27</intersection>
<intersection>120 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>101,45,101,45.5</points>
<connection>
<GID>547</GID>
<name>N_in1</name></connection>
<intersection>45 2</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>117,49.5,117,52</points>
<connection>
<GID>552</GID>
<name>IN_0</name></connection>
<intersection>49.5 14</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>113.5,70,120,70</points>
<intersection>113.5 32</intersection>
<intersection>120 0</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>113.5,70,113.5,72</points>
<connection>
<GID>541</GID>
<name>IN_0</name></connection>
<intersection>70 30</intersection></vsegment></shape></wire>
<wire>
<ID>453</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>111,67.5,113,67.5</points>
<connection>
<GID>542</GID>
<name>OUT</name></connection>
<connection>
<GID>540</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>454</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,44.5,102,76</points>
<connection>
<GID>546</GID>
<name>N_in0</name></connection>
<connection>
<GID>545</GID>
<name>N_in1</name></connection>
<intersection>44.5 6</intersection>
<intersection>66.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>102,66.5,105,66.5</points>
<connection>
<GID>542</GID>
<name>IN_1</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>102,44.5,124.5,44.5</points>
<intersection>102 0</intersection>
<intersection>124.5 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>124.5,44.5,124.5,50.5</points>
<connection>
<GID>560</GID>
<name>IN_0</name></connection>
<intersection>44.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>455</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,72.5,108,74</points>
<connection>
<GID>542</GID>
<name>SEL_1</name></connection>
<intersection>74 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,74,123,74</points>
<connection>
<GID>553</GID>
<name>N_in0</name></connection>
<connection>
<GID>549</GID>
<name>N_in1</name></connection>
<intersection>108 0</intersection></hsegment></shape></wire>
<wire>
<ID>456</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109,72.5,109,75</points>
<connection>
<GID>542</GID>
<name>SEL_0</name></connection>
<intersection>75 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,75,123,75</points>
<connection>
<GID>554</GID>
<name>N_in0</name></connection>
<connection>
<GID>550</GID>
<name>N_in1</name></connection>
<intersection>109 0</intersection></hsegment></shape></wire>
<wire>
<ID>457</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,62.5,113,64.5</points>
<connection>
<GID>540</GID>
<name>clock</name></connection>
<intersection>62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111.5,62.5,113,62.5</points>
<connection>
<GID>556</GID>
<name>IN_0</name></connection>
<intersection>113 0</intersection></hsegment></shape></wire>
<wire>
<ID>458</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,60.5,116,61.5</points>
<connection>
<GID>540</GID>
<name>clear</name></connection>
<intersection>60.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>111.5,60.5,116,60.5</points>
<connection>
<GID>558</GID>
<name>IN_0</name></connection>
<intersection>116 0</intersection></hsegment></shape></wire>
<wire>
<ID>459</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,55,110,57.5</points>
<intersection>55 1</intersection>
<intersection>57.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109.5,55,110,55</points>
<connection>
<GID>557</GID>
<name>IN_2</name></connection>
<intersection>110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,57.5,111,57.5</points>
<connection>
<GID>551</GID>
<name>OUT</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>460</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109.5,53,111,53</points>
<connection>
<GID>557</GID>
<name>IN_1</name></connection>
<connection>
<GID>552</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>461</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,48.5,110,51</points>
<intersection>48.5 1</intersection>
<intersection>51 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110,48.5,111,48.5</points>
<connection>
<GID>555</GID>
<name>OUT</name></connection>
<intersection>110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109.5,51,110,51</points>
<connection>
<GID>557</GID>
<name>IN_0</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>462</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>98.5,53,103.5,53</points>
<connection>
<GID>559</GID>
<name>N_in1</name></connection>
<connection>
<GID>557</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>463</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,53,121,58.5</points>
<intersection>53 8</intersection>
<intersection>54 1</intersection>
<intersection>58.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117,54,121,54</points>
<connection>
<GID>552</GID>
<name>IN_1</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>117,58.5,121,58.5</points>
<connection>
<GID>551</GID>
<name>IN_1</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>121,53,123,53</points>
<connection>
<GID>539</GID>
<name>N_in0</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>464</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,47.5,119,56.5</points>
<intersection>47.5 3</intersection>
<intersection>50.5 2</intersection>
<intersection>56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117,56.5,119,56.5</points>
<connection>
<GID>551</GID>
<name>IN_0</name></connection>
<intersection>119 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>119,50.5,120.5,50.5</points>
<connection>
<GID>560</GID>
<name>OUT_0</name></connection>
<intersection>119 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>117,47.5,119,47.5</points>
<connection>
<GID>555</GID>
<name>IN_0</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>465</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,45.5,99.5,70.5</points>
<intersection>45.5 2</intersection>
<intersection>70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99.5,70.5,105,70.5</points>
<connection>
<GID>542</GID>
<name>IN_3</name></connection>
<intersection>99.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99.5,45.5,100,45.5</points>
<connection>
<GID>544</GID>
<name>N_in1</name></connection>
<intersection>99.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>466</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,68.5,101,76</points>
<connection>
<GID>548</GID>
<name>N_in0</name></connection>
<intersection>68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,68.5,105,68.5</points>
<connection>
<GID>542</GID>
<name>IN_2</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>467</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,53,96.5,53</points>
<connection>
<GID>559</GID>
<name>N_in0</name></connection>
<connection>
<GID>613</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>468</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,75,96.5,75</points>
<connection>
<GID>550</GID>
<name>N_in0</name></connection>
<connection>
<GID>608</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>469</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,74,96.5,74</points>
<connection>
<GID>549</GID>
<name>N_in0</name></connection>
<connection>
<GID>610</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>470</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148.5,45,148.5,70</points>
<intersection>45 2</intersection>
<intersection>49.5 14</intersection>
<intersection>67.5 7</intersection>
<intersection>70 30</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>128.5,45,148.5,45</points>
<intersection>128.5 4</intersection>
<intersection>129.5 17</intersection>
<intersection>148.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>128.5,45,128.5,76</points>
<connection>
<GID>565</GID>
<name>N_in0</name></connection>
<intersection>45 2</intersection>
<intersection>64.5 9</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>147.5,67.5,148.5,67.5</points>
<connection>
<GID>562</GID>
<name>OUT_0</name></connection>
<intersection>148.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>128.5,64.5,133.5,64.5</points>
<connection>
<GID>564</GID>
<name>IN_0</name></connection>
<intersection>128.5 4</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>145.5,49.5,148.5,49.5</points>
<connection>
<GID>577</GID>
<name>IN_1</name></connection>
<intersection>145.5 27</intersection>
<intersection>148.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>129.5,45,129.5,45.5</points>
<connection>
<GID>569</GID>
<name>N_in1</name></connection>
<intersection>45 2</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>145.5,49.5,145.5,52</points>
<connection>
<GID>574</GID>
<name>IN_0</name></connection>
<intersection>49.5 14</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>142,70,148.5,70</points>
<intersection>142 32</intersection>
<intersection>148.5 0</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>142,70,142,72</points>
<connection>
<GID>563</GID>
<name>IN_0</name></connection>
<intersection>70 30</intersection></vsegment></shape></wire>
<wire>
<ID>471</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>139.5,67.5,141.5,67.5</points>
<connection>
<GID>564</GID>
<name>OUT</name></connection>
<connection>
<GID>562</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>472</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,44.5,130.5,76</points>
<connection>
<GID>568</GID>
<name>N_in0</name></connection>
<connection>
<GID>567</GID>
<name>N_in1</name></connection>
<intersection>44.5 6</intersection>
<intersection>66.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>130.5,66.5,133.5,66.5</points>
<connection>
<GID>564</GID>
<name>IN_1</name></connection>
<intersection>130.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>130.5,44.5,153,44.5</points>
<intersection>130.5 0</intersection>
<intersection>153 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>153,44.5,153,50.5</points>
<connection>
<GID>583</GID>
<name>IN_0</name></connection>
<intersection>44.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>473</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136.5,72.5,136.5,74</points>
<connection>
<GID>564</GID>
<name>SEL_1</name></connection>
<intersection>74 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,74,151.5,74</points>
<connection>
<GID>575</GID>
<name>N_in0</name></connection>
<connection>
<GID>571</GID>
<name>N_in1</name></connection>
<intersection>136.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>474</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137.5,72.5,137.5,75</points>
<connection>
<GID>564</GID>
<name>SEL_0</name></connection>
<intersection>75 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,75,151.5,75</points>
<connection>
<GID>576</GID>
<name>N_in0</name></connection>
<connection>
<GID>572</GID>
<name>N_in1</name></connection>
<intersection>137.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>475</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,62.5,141.5,64.5</points>
<connection>
<GID>562</GID>
<name>clock</name></connection>
<intersection>62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>140,62.5,141.5,62.5</points>
<connection>
<GID>578</GID>
<name>IN_0</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>476</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144.5,60.5,144.5,61.5</points>
<connection>
<GID>562</GID>
<name>clear</name></connection>
<intersection>60.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>140,60.5,144.5,60.5</points>
<connection>
<GID>580</GID>
<name>IN_0</name></connection>
<intersection>144.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>477</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,55,138.5,57.5</points>
<intersection>55 1</intersection>
<intersection>57.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,55,138.5,55</points>
<connection>
<GID>579</GID>
<name>IN_2</name></connection>
<intersection>138.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138.5,57.5,139.5,57.5</points>
<connection>
<GID>573</GID>
<name>OUT</name></connection>
<intersection>138.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>478</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>138,53,139.5,53</points>
<connection>
<GID>579</GID>
<name>IN_1</name></connection>
<connection>
<GID>574</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>479</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,48.5,138.5,51</points>
<intersection>48.5 1</intersection>
<intersection>51 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138.5,48.5,139.5,48.5</points>
<connection>
<GID>577</GID>
<name>OUT</name></connection>
<intersection>138.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138,51,138.5,51</points>
<connection>
<GID>579</GID>
<name>IN_0</name></connection>
<intersection>138.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>480</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>127,53,132,53</points>
<connection>
<GID>581</GID>
<name>N_in1</name></connection>
<connection>
<GID>579</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>481</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149.5,53,149.5,58.5</points>
<intersection>53 8</intersection>
<intersection>54 1</intersection>
<intersection>58.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145.5,54,149.5,54</points>
<connection>
<GID>574</GID>
<name>IN_1</name></connection>
<intersection>149.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>145.5,58.5,149.5,58.5</points>
<connection>
<GID>573</GID>
<name>IN_1</name></connection>
<intersection>149.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>149.5,53,151.5,53</points>
<connection>
<GID>561</GID>
<name>N_in0</name></connection>
<intersection>149.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>482</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147.5,47.5,147.5,56.5</points>
<intersection>47.5 3</intersection>
<intersection>50.5 2</intersection>
<intersection>56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145.5,56.5,147.5,56.5</points>
<connection>
<GID>573</GID>
<name>IN_0</name></connection>
<intersection>147.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>147.5,50.5,149,50.5</points>
<connection>
<GID>583</GID>
<name>OUT_0</name></connection>
<intersection>147.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>145.5,47.5,147.5,47.5</points>
<connection>
<GID>577</GID>
<name>IN_0</name></connection>
<intersection>147.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>483</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,45.5,128,70.5</points>
<intersection>45.5 2</intersection>
<intersection>70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128,70.5,133.5,70.5</points>
<connection>
<GID>564</GID>
<name>IN_3</name></connection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>128,45.5,128.5,45.5</points>
<connection>
<GID>566</GID>
<name>N_in1</name></connection>
<intersection>128 0</intersection></hsegment></shape></wire>
<wire>
<ID>506</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,68.5,129.5,76</points>
<connection>
<GID>570</GID>
<name>N_in0</name></connection>
<intersection>68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,68.5,133.5,68.5</points>
<connection>
<GID>564</GID>
<name>IN_2</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>507</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,75,125,75</points>
<connection>
<GID>554</GID>
<name>N_in1</name></connection>
<connection>
<GID>572</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>508</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,74,125,74</points>
<connection>
<GID>553</GID>
<name>N_in1</name></connection>
<connection>
<GID>571</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>509</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,53,125,53</points>
<connection>
<GID>539</GID>
<name>N_in1</name></connection>
<connection>
<GID>581</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>510</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177,45,177,70</points>
<intersection>45 2</intersection>
<intersection>49.5 14</intersection>
<intersection>67.5 7</intersection>
<intersection>70 30</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>157,45,177,45</points>
<intersection>157 4</intersection>
<intersection>158 17</intersection>
<intersection>177 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>157,45,157,76</points>
<connection>
<GID>589</GID>
<name>N_in0</name></connection>
<intersection>45 2</intersection>
<intersection>64.5 9</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>176,67.5,177,67.5</points>
<connection>
<GID>586</GID>
<name>OUT_0</name></connection>
<intersection>177 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>157,64.5,162,64.5</points>
<connection>
<GID>588</GID>
<name>IN_0</name></connection>
<intersection>157 4</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>174,49.5,177,49.5</points>
<connection>
<GID>601</GID>
<name>IN_1</name></connection>
<intersection>174 27</intersection>
<intersection>177 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>158,45,158,45.5</points>
<connection>
<GID>593</GID>
<name>N_in1</name></connection>
<intersection>45 2</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>174,49.5,174,52</points>
<connection>
<GID>598</GID>
<name>IN_0</name></connection>
<intersection>49.5 14</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>170.5,70,177,70</points>
<intersection>170.5 32</intersection>
<intersection>177 0</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>170.5,70,170.5,72</points>
<connection>
<GID>587</GID>
<name>IN_0</name></connection>
<intersection>70 30</intersection></vsegment></shape></wire>
<wire>
<ID>511</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>168,67.5,170,67.5</points>
<connection>
<GID>588</GID>
<name>OUT</name></connection>
<connection>
<GID>586</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>512</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,44.5,159,76</points>
<connection>
<GID>592</GID>
<name>N_in0</name></connection>
<connection>
<GID>591</GID>
<name>N_in1</name></connection>
<intersection>44.5 6</intersection>
<intersection>66.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>159,66.5,162,66.5</points>
<connection>
<GID>588</GID>
<name>IN_1</name></connection>
<intersection>159 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>159,44.5,181.5,44.5</points>
<intersection>159 0</intersection>
<intersection>181.5 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>181.5,44.5,181.5,50.5</points>
<connection>
<GID>612</GID>
<name>IN_0</name></connection>
<intersection>44.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>513</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165,72.5,165,74</points>
<connection>
<GID>588</GID>
<name>SEL_1</name></connection>
<intersection>74 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>155.5,74,180,74</points>
<connection>
<GID>599</GID>
<name>N_in0</name></connection>
<connection>
<GID>595</GID>
<name>N_in1</name></connection>
<intersection>165 0</intersection></hsegment></shape></wire>
<wire>
<ID>514</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,72.5,166,75</points>
<connection>
<GID>588</GID>
<name>SEL_0</name></connection>
<intersection>75 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>155.5,75,180,75</points>
<connection>
<GID>600</GID>
<name>N_in0</name></connection>
<connection>
<GID>596</GID>
<name>N_in1</name></connection>
<intersection>166 0</intersection></hsegment></shape></wire>
<wire>
<ID>515</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,62.5,170,64.5</points>
<connection>
<GID>586</GID>
<name>clock</name></connection>
<intersection>62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168.5,62.5,170,62.5</points>
<connection>
<GID>602</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment></shape></wire>
<wire>
<ID>516</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173,60.5,173,61.5</points>
<connection>
<GID>586</GID>
<name>clear</name></connection>
<intersection>60.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>168.5,60.5,173,60.5</points>
<connection>
<GID>607</GID>
<name>IN_0</name></connection>
<intersection>173 0</intersection></hsegment></shape></wire>
<wire>
<ID>517</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,55,167,57.5</points>
<intersection>55 1</intersection>
<intersection>57.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166.5,55,167,55</points>
<connection>
<GID>604</GID>
<name>IN_2</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>167,57.5,168,57.5</points>
<connection>
<GID>597</GID>
<name>OUT</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>518</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>166.5,53,168,53</points>
<connection>
<GID>604</GID>
<name>IN_1</name></connection>
<connection>
<GID>598</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>519</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,48.5,167,51</points>
<intersection>48.5 1</intersection>
<intersection>51 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167,48.5,168,48.5</points>
<connection>
<GID>601</GID>
<name>OUT</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>166.5,51,167,51</points>
<connection>
<GID>604</GID>
<name>IN_0</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>520</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>155.5,53,160.5,53</points>
<connection>
<GID>609</GID>
<name>N_in1</name></connection>
<connection>
<GID>604</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>521</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178,53,178,58.5</points>
<intersection>53 8</intersection>
<intersection>54 1</intersection>
<intersection>58.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>174,54,178,54</points>
<connection>
<GID>598</GID>
<name>IN_1</name></connection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>174,58.5,178,58.5</points>
<connection>
<GID>597</GID>
<name>IN_1</name></connection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>178,53,180,53</points>
<connection>
<GID>584</GID>
<name>N_in0</name></connection>
<intersection>178 0</intersection></hsegment></shape></wire>
<wire>
<ID>522</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176,47.5,176,56.5</points>
<intersection>47.5 3</intersection>
<intersection>50.5 2</intersection>
<intersection>56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>174,56.5,176,56.5</points>
<connection>
<GID>597</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>176,50.5,177.5,50.5</points>
<connection>
<GID>612</GID>
<name>OUT_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>174,47.5,176,47.5</points>
<connection>
<GID>601</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment></shape></wire>
<wire>
<ID>523</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,45.5,156.5,70.5</points>
<intersection>45.5 2</intersection>
<intersection>70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156.5,70.5,162,70.5</points>
<connection>
<GID>588</GID>
<name>IN_3</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156.5,45.5,157,45.5</points>
<connection>
<GID>590</GID>
<name>N_in1</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>524</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158,68.5,158,76</points>
<connection>
<GID>594</GID>
<name>N_in0</name></connection>
<intersection>68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>158,68.5,162,68.5</points>
<connection>
<GID>588</GID>
<name>IN_2</name></connection>
<intersection>158 0</intersection></hsegment></shape></wire>
<wire>
<ID>525</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153.5,53,153.5,53</points>
<connection>
<GID>561</GID>
<name>N_in1</name></connection>
<connection>
<GID>609</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>526</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153.5,75,153.5,75</points>
<connection>
<GID>576</GID>
<name>N_in1</name></connection>
<connection>
<GID>596</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>527</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153.5,74,153.5,74</points>
<connection>
<GID>575</GID>
<name>N_in1</name></connection>
<connection>
<GID>595</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>528</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205.5,45,205.5,70</points>
<intersection>45 2</intersection>
<intersection>49.5 14</intersection>
<intersection>67.5 7</intersection>
<intersection>70 30</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>185.5,45,205.5,45</points>
<intersection>185.5 4</intersection>
<intersection>186.5 17</intersection>
<intersection>205.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>185.5,45,185.5,76</points>
<connection>
<GID>620</GID>
<name>N_in0</name></connection>
<intersection>45 2</intersection>
<intersection>64.5 9</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>204.5,67.5,205.5,67.5</points>
<connection>
<GID>616</GID>
<name>OUT_0</name></connection>
<intersection>205.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>185.5,64.5,190.5,64.5</points>
<connection>
<GID>619</GID>
<name>IN_0</name></connection>
<intersection>185.5 4</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>202.5,49.5,205.5,49.5</points>
<connection>
<GID>530</GID>
<name>IN_1</name></connection>
<intersection>202.5 27</intersection>
<intersection>205.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>186.5,45,186.5,45.5</points>
<connection>
<GID>520</GID>
<name>N_in1</name></connection>
<intersection>45 2</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>202.5,49.5,202.5,52</points>
<connection>
<GID>527</GID>
<name>IN_0</name></connection>
<intersection>49.5 14</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>199,70,205.5,70</points>
<intersection>199 32</intersection>
<intersection>205.5 0</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>199,70,199,72</points>
<connection>
<GID>618</GID>
<name>IN_0</name></connection>
<intersection>70 30</intersection></vsegment></shape></wire>
<wire>
<ID>529</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>196.5,67.5,198.5,67.5</points>
<connection>
<GID>619</GID>
<name>OUT</name></connection>
<connection>
<GID>616</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>530</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,44.5,187.5,76</points>
<connection>
<GID>625</GID>
<name>N_in0</name></connection>
<connection>
<GID>622</GID>
<name>N_in1</name></connection>
<intersection>44.5 6</intersection>
<intersection>66.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>187.5,66.5,190.5,66.5</points>
<connection>
<GID>619</GID>
<name>IN_1</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>187.5,44.5,210,44.5</points>
<intersection>187.5 0</intersection>
<intersection>210 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>210,44.5,210,50.5</points>
<connection>
<GID>535</GID>
<name>IN_0</name></connection>
<intersection>44.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>531</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>193.5,72.5,193.5,74</points>
<connection>
<GID>619</GID>
<name>SEL_1</name></connection>
<intersection>74 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184,74,208.5,74</points>
<connection>
<GID>528</GID>
<name>N_in0</name></connection>
<connection>
<GID>524</GID>
<name>N_in1</name></connection>
<intersection>193.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>532</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,72.5,194.5,75</points>
<connection>
<GID>619</GID>
<name>SEL_0</name></connection>
<intersection>75 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184,75,208.5,75</points>
<connection>
<GID>529</GID>
<name>N_in0</name></connection>
<connection>
<GID>525</GID>
<name>N_in1</name></connection>
<intersection>194.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>533</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,62.5,198.5,64.5</points>
<connection>
<GID>616</GID>
<name>clock</name></connection>
<intersection>62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>197,62.5,198.5,62.5</points>
<connection>
<GID>531</GID>
<name>IN_0</name></connection>
<intersection>198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>534</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201.5,60.5,201.5,61.5</points>
<connection>
<GID>616</GID>
<name>clear</name></connection>
<intersection>60.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>197,60.5,201.5,60.5</points>
<connection>
<GID>533</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>535</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>195.5,55,195.5,57.5</points>
<intersection>55 1</intersection>
<intersection>57.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>195,55,195.5,55</points>
<connection>
<GID>532</GID>
<name>IN_2</name></connection>
<intersection>195.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>195.5,57.5,196.5,57.5</points>
<connection>
<GID>526</GID>
<name>OUT</name></connection>
<intersection>195.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>536</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,53,196.5,53</points>
<connection>
<GID>532</GID>
<name>IN_1</name></connection>
<connection>
<GID>527</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>537</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>195.5,48.5,195.5,51</points>
<intersection>48.5 1</intersection>
<intersection>51 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>195.5,48.5,196.5,48.5</points>
<connection>
<GID>530</GID>
<name>OUT</name></connection>
<intersection>195.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>195,51,195.5,51</points>
<connection>
<GID>532</GID>
<name>IN_0</name></connection>
<intersection>195.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>538</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>184,53,189,53</points>
<connection>
<GID>534</GID>
<name>N_in1</name></connection>
<connection>
<GID>532</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>539</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206.5,53,206.5,58.5</points>
<intersection>53 8</intersection>
<intersection>54 1</intersection>
<intersection>58.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>202.5,54,206.5,54</points>
<connection>
<GID>527</GID>
<name>IN_1</name></connection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>202.5,58.5,206.5,58.5</points>
<connection>
<GID>526</GID>
<name>IN_1</name></connection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>206.5,53,208.5,53</points>
<connection>
<GID>614</GID>
<name>N_in0</name></connection>
<intersection>206.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>540</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204.5,47.5,204.5,56.5</points>
<intersection>47.5 3</intersection>
<intersection>50.5 2</intersection>
<intersection>56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>202.5,56.5,204.5,56.5</points>
<connection>
<GID>526</GID>
<name>IN_0</name></connection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>204.5,50.5,206,50.5</points>
<connection>
<GID>535</GID>
<name>OUT_0</name></connection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>202.5,47.5,204.5,47.5</points>
<connection>
<GID>530</GID>
<name>IN_0</name></connection>
<intersection>204.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>541</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,45.5,185,70.5</points>
<intersection>45.5 2</intersection>
<intersection>70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185,70.5,190.5,70.5</points>
<connection>
<GID>619</GID>
<name>IN_3</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>185,45.5,185.5,45.5</points>
<connection>
<GID>621</GID>
<name>N_in1</name></connection>
<intersection>185 0</intersection></hsegment></shape></wire>
<wire>
<ID>542</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186.5,68.5,186.5,76</points>
<connection>
<GID>522</GID>
<name>N_in0</name></connection>
<intersection>68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>186.5,68.5,190.5,68.5</points>
<connection>
<GID>619</GID>
<name>IN_2</name></connection>
<intersection>186.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>543</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182,53,182,53</points>
<connection>
<GID>534</GID>
<name>N_in0</name></connection>
<connection>
<GID>584</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>544</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182,75,182,75</points>
<connection>
<GID>525</GID>
<name>N_in0</name></connection>
<connection>
<GID>600</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>545</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182,74,182,74</points>
<connection>
<GID>524</GID>
<name>N_in0</name></connection>
<connection>
<GID>599</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>546</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210.5,53,210.5,53</points>
<connection>
<GID>537</GID>
<name>N_in0</name></connection>
<connection>
<GID>614</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>547</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211.5,54,211.5,76</points>
<connection>
<GID>537</GID>
<name>N_in3</name></connection>
<connection>
<GID>536</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>548</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211.5,45.5,211.5,52</points>
<connection>
<GID>538</GID>
<name>N_in1</name></connection>
<connection>
<GID>537</GID>
<name>N_in2</name></connection></vsegment></shape></wire>
<wire>
<ID>549</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,45.5,80,76</points>
<connection>
<GID>617</GID>
<name>N_in1</name></connection>
<connection>
<GID>615</GID>
<name>N_in0</name></connection>
<intersection>68.5 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>80,68.5,81.5,68.5</points>
<connection>
<GID>523</GID>
<name>IN_0</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>550</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>80.5,53,94.5,53</points>
<connection>
<GID>613</GID>
<name>N_in0</name></connection>
<intersection>80.5 8</intersection>
<intersection>81 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>81,45.5,81,53</points>
<connection>
<GID>605</GID>
<name>N_in1</name></connection>
<intersection>53 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>80.5,53,80.5,71</points>
<intersection>53 2</intersection>
<intersection>71 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>80.5,71,81.5,71</points>
<connection>
<GID>624</GID>
<name>IN_1</name></connection>
<intersection>80.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>551</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,70.5,87.5,72</points>
<connection>
<GID>626</GID>
<name>IN_0</name></connection>
<connection>
<GID>624</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>552</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,69.5,93.5,75</points>
<connection>
<GID>626</GID>
<name>OUT</name></connection>
<intersection>75 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93.5,75,94.5,75</points>
<connection>
<GID>608</GID>
<name>N_in0</name></connection>
<intersection>93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>553</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94.5,64.5,94.5,74</points>
<connection>
<GID>610</GID>
<name>N_in0</name></connection>
<intersection>64.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>93.5,64.5,94.5,64.5</points>
<connection>
<GID>521</GID>
<name>OUT</name></connection>
<intersection>94.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>554</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,63.5,81,76</points>
<connection>
<GID>603</GID>
<name>N_in0</name></connection>
<intersection>63.5 3</intersection>
<intersection>73 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81,73,81.5,73</points>
<connection>
<GID>624</GID>
<name>IN_0</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>81,63.5,87.5,63.5</points>
<connection>
<GID>521</GID>
<name>IN_1</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>555</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,68.5,87.5,68.5</points>
<connection>
<GID>626</GID>
<name>IN_1</name></connection>
<connection>
<GID>523</GID>
<name>OUT_0</name></connection>
<intersection>86.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>86.5,65.5,86.5,68.5</points>
<intersection>65.5 8</intersection>
<intersection>68.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>86.5,65.5,87.5,65.5</points>
<connection>
<GID>521</GID>
<name>IN_0</name></connection>
<intersection>86.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>556</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211.5,78,211.5,78</points>
<connection>
<GID>436</GID>
<name>N_in0</name></connection>
<connection>
<GID>536</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>557</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186.5,78,186.5,78</points>
<connection>
<GID>418</GID>
<name>N_in0</name></connection>
<connection>
<GID>522</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>558</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,78,100,78</points>
<connection>
<GID>442</GID>
<name>N_in0</name></connection>
<connection>
<GID>543</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>559</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128.5,78,128.5,78</points>
<connection>
<GID>464</GID>
<name>N_in0</name></connection>
<connection>
<GID>565</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>560</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,78,102,78</points>
<connection>
<GID>443</GID>
<name>N_in0</name></connection>
<connection>
<GID>546</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>561</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,78,101,78</points>
<connection>
<GID>445</GID>
<name>N_in0</name></connection>
<connection>
<GID>548</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>562</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,78,130.5,78</points>
<connection>
<GID>465</GID>
<name>N_in0</name></connection>
<connection>
<GID>568</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>563</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,78,129.5,78</points>
<connection>
<GID>467</GID>
<name>N_in0</name></connection>
<connection>
<GID>570</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>564</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157,78,157,78</points>
<connection>
<GID>486</GID>
<name>N_in0</name></connection>
<connection>
<GID>589</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>565</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,78,159,78</points>
<connection>
<GID>487</GID>
<name>N_in0</name></connection>
<connection>
<GID>592</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,148.5,120,173.5</points>
<intersection>148.5 2</intersection>
<intersection>153 14</intersection>
<intersection>171 7</intersection>
<intersection>173.5 30</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>100,148.5,120,148.5</points>
<intersection>100 4</intersection>
<intersection>101 17</intersection>
<intersection>120 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>100,148.5,100,179.5</points>
<connection>
<GID>236</GID>
<name>N_in0</name></connection>
<intersection>148.5 2</intersection>
<intersection>168 9</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>119,171,120,171</points>
<connection>
<GID>233</GID>
<name>OUT_0</name></connection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>100,168,105,168</points>
<connection>
<GID>235</GID>
<name>IN_0</name></connection>
<intersection>100 4</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>117,153,120,153</points>
<connection>
<GID>248</GID>
<name>IN_1</name></connection>
<intersection>117 27</intersection>
<intersection>120 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>101,148.5,101,149</points>
<connection>
<GID>240</GID>
<name>N_in1</name></connection>
<intersection>148.5 2</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>117,153,117,155.5</points>
<connection>
<GID>245</GID>
<name>IN_0</name></connection>
<intersection>153 14</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>113.5,173.5,120,173.5</points>
<intersection>113.5 32</intersection>
<intersection>120 0</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>113.5,173.5,113.5,175.5</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<intersection>173.5 30</intersection></vsegment></shape></wire>
<wire>
<ID>566</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158,78,158,78</points>
<connection>
<GID>489</GID>
<name>N_in0</name></connection>
<connection>
<GID>594</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>111,171,113,171</points>
<connection>
<GID>235</GID>
<name>OUT</name></connection>
<connection>
<GID>233</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>567</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,78,81,78</points>
<connection>
<GID>501</GID>
<name>N_in0</name></connection>
<connection>
<GID>603</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,148,102,179.5</points>
<connection>
<GID>238</GID>
<name>N_in1</name></connection>
<connection>
<GID>239</GID>
<name>N_in0</name></connection>
<intersection>148 6</intersection>
<intersection>170 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>102,170,105,170</points>
<connection>
<GID>235</GID>
<name>IN_1</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>102,148,124.5,148</points>
<intersection>102 0</intersection>
<intersection>124.5 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>124.5,148,124.5,154</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<intersection>148 6</intersection></vsegment></shape></wire>
<wire>
<ID>568</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,78,80,78</points>
<connection>
<GID>511</GID>
<name>N_in0</name></connection>
<connection>
<GID>615</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,176,108,177.5</points>
<connection>
<GID>235</GID>
<name>SEL_1</name></connection>
<intersection>177.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,177.5,123,177.5</points>
<connection>
<GID>242</GID>
<name>N_in1</name></connection>
<connection>
<GID>246</GID>
<name>N_in0</name></connection>
<intersection>108 0</intersection></hsegment></shape></wire>
<wire>
<ID>569</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185.5,78,185.5,78</points>
<connection>
<GID>515</GID>
<name>N_in0</name></connection>
<connection>
<GID>620</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109,176,109,178.5</points>
<connection>
<GID>235</GID>
<name>SEL_0</name></connection>
<intersection>178.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,178.5,123,178.5</points>
<connection>
<GID>243</GID>
<name>N_in1</name></connection>
<connection>
<GID>247</GID>
<name>N_in0</name></connection>
<intersection>109 0</intersection></hsegment></shape></wire>
<wire>
<ID>570</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,78,187.5,78</points>
<connection>
<GID>516</GID>
<name>N_in0</name></connection>
<connection>
<GID>625</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,166,113,168</points>
<connection>
<GID>233</GID>
<name>clock</name></connection>
<intersection>166 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111.5,166,113,166</points>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<intersection>113 0</intersection></hsegment></shape></wire>
<wire>
<ID>571</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,181.5,81,182.5</points>
<connection>
<GID>295</GID>
<name>N_in1</name></connection>
<connection>
<GID>628</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,164,116,165</points>
<connection>
<GID>233</GID>
<name>clear</name></connection>
<intersection>164 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>111.5,164,116,164</points>
<connection>
<GID>251</GID>
<name>IN_0</name></connection>
<intersection>116 0</intersection></hsegment></shape></wire>
<wire>
<ID>572</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,42,80,43.5</points>
<connection>
<GID>617</GID>
<name>N_in0</name></connection>
<intersection>42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79,42,80,42</points>
<connection>
<GID>633</GID>
<name>IN_0</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,158.5,110,161</points>
<intersection>158.5 1</intersection>
<intersection>161 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109.5,158.5,110,158.5</points>
<connection>
<GID>250</GID>
<name>IN_2</name></connection>
<intersection>110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,161,111,161</points>
<connection>
<GID>244</GID>
<name>OUT</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>573</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211.5,42.5,211.5,43.5</points>
<connection>
<GID>538</GID>
<name>N_in0</name></connection>
<connection>
<GID>635</GID>
<name>OUT_0</name></connection>
<intersection>42.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>100,42.5,211.5,42.5</points>
<intersection>100 11</intersection>
<intersection>128.5 9</intersection>
<intersection>157 6</intersection>
<intersection>185.5 7</intersection>
<intersection>211.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>157,42.5,157,43.5</points>
<connection>
<GID>590</GID>
<name>N_in0</name></connection>
<intersection>42.5 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>185.5,42.5,185.5,43.5</points>
<connection>
<GID>621</GID>
<name>N_in0</name></connection>
<intersection>42.5 4</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>128.5,42.5,128.5,43.5</points>
<connection>
<GID>566</GID>
<name>N_in0</name></connection>
<intersection>42.5 4</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>100,42.5,100,43.5</points>
<connection>
<GID>544</GID>
<name>N_in0</name></connection>
<intersection>42.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109.5,156.5,111,156.5</points>
<connection>
<GID>250</GID>
<name>IN_1</name></connection>
<connection>
<GID>245</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>574</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101,182.5,211.5,182.5</points>
<intersection>101 10</intersection>
<intersection>129.5 8</intersection>
<intersection>158 6</intersection>
<intersection>186.5 3</intersection>
<intersection>211.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>186.5,181.5,186.5,182.5</points>
<connection>
<GID>215</GID>
<name>N_in1</name></connection>
<intersection>182.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>211.5,181.5,211.5,182.5</points>
<connection>
<GID>229</GID>
<name>N_in1</name></connection>
<intersection>182.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>158,181.5,158,182.5</points>
<connection>
<GID>286</GID>
<name>N_in1</name></connection>
<intersection>182.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>129.5,181.5,129.5,182.5</points>
<connection>
<GID>263</GID>
<name>N_in1</name></connection>
<intersection>182.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>101,181.5,101,182.5</points>
<connection>
<GID>241</GID>
<name>N_in1</name></connection>
<intersection>182.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,152,110,154.5</points>
<intersection>152 1</intersection>
<intersection>154.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110,152,111,152</points>
<connection>
<GID>248</GID>
<name>OUT</name></connection>
<intersection>110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109.5,154.5,110,154.5</points>
<connection>
<GID>250</GID>
<name>IN_0</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>575</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,39,102,43.5</points>
<connection>
<GID>545</GID>
<name>N_in0</name></connection>
<intersection>39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,39,102,39</points>
<connection>
<GID>636</GID>
<name>IN_0</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>98.5,156.5,103.5,156.5</points>
<connection>
<GID>252</GID>
<name>N_in1</name></connection>
<connection>
<GID>250</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>576</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,37,130.5,43.5</points>
<connection>
<GID>567</GID>
<name>N_in0</name></connection>
<intersection>37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,37,130.5,37</points>
<connection>
<GID>638</GID>
<name>IN_0</name></connection>
<intersection>130.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,156.5,121,162</points>
<intersection>156.5 8</intersection>
<intersection>157.5 1</intersection>
<intersection>162 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117,157.5,121,157.5</points>
<connection>
<GID>245</GID>
<name>IN_1</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>117,162,121,162</points>
<connection>
<GID>244</GID>
<name>IN_1</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>121,156.5,123,156.5</points>
<connection>
<GID>232</GID>
<name>N_in0</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>577</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,35,159,43.5</points>
<connection>
<GID>591</GID>
<name>N_in0</name></connection>
<intersection>35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,35,159,35</points>
<connection>
<GID>639</GID>
<name>IN_0</name></connection>
<intersection>159 0</intersection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,151,119,160</points>
<intersection>151 3</intersection>
<intersection>154 2</intersection>
<intersection>160 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117,160,119,160</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<intersection>119 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>119,154,120.5,154</points>
<connection>
<GID>253</GID>
<name>OUT_0</name></connection>
<intersection>119 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>117,151,119,151</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>578</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,33,187.5,43.5</points>
<connection>
<GID>622</GID>
<name>N_in0</name></connection>
<intersection>33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,33,187.5,33</points>
<connection>
<GID>640</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,149,99.5,174</points>
<intersection>149 2</intersection>
<intersection>174 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99.5,174,105,174</points>
<connection>
<GID>235</GID>
<name>IN_3</name></connection>
<intersection>99.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99.5,149,100,149</points>
<connection>
<GID>237</GID>
<name>N_in1</name></connection>
<intersection>99.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,172,101,179.5</points>
<connection>
<GID>241</GID>
<name>N_in0</name></connection>
<intersection>172 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,172,105,172</points>
<connection>
<GID>235</GID>
<name>IN_2</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,156.5,96.5,156.5</points>
<connection>
<GID>252</GID>
<name>N_in0</name></connection>
<connection>
<GID>303</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,178.5,96.5,178.5</points>
<connection>
<GID>243</GID>
<name>N_in0</name></connection>
<connection>
<GID>299</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,177.5,96.5,177.5</points>
<connection>
<GID>242</GID>
<name>N_in0</name></connection>
<connection>
<GID>301</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148.5,148.5,148.5,173.5</points>
<intersection>148.5 2</intersection>
<intersection>153 14</intersection>
<intersection>171 7</intersection>
<intersection>173.5 30</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>128.5,148.5,148.5,148.5</points>
<intersection>128.5 4</intersection>
<intersection>129.5 17</intersection>
<intersection>148.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>128.5,148.5,128.5,179.5</points>
<connection>
<GID>258</GID>
<name>N_in0</name></connection>
<intersection>148.5 2</intersection>
<intersection>168 9</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>147.5,171,148.5,171</points>
<connection>
<GID>255</GID>
<name>OUT_0</name></connection>
<intersection>148.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>128.5,168,133.5,168</points>
<connection>
<GID>257</GID>
<name>IN_0</name></connection>
<intersection>128.5 4</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>145.5,153,148.5,153</points>
<connection>
<GID>270</GID>
<name>IN_1</name></connection>
<intersection>145.5 27</intersection>
<intersection>148.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>129.5,148.5,129.5,149</points>
<connection>
<GID>262</GID>
<name>N_in1</name></connection>
<intersection>148.5 2</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>145.5,153,145.5,155.5</points>
<connection>
<GID>267</GID>
<name>IN_0</name></connection>
<intersection>153 14</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>142,173.5,148.5,173.5</points>
<intersection>142 32</intersection>
<intersection>148.5 0</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>142,173.5,142,175.5</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<intersection>173.5 30</intersection></vsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>139.5,171,141.5,171</points>
<connection>
<GID>257</GID>
<name>OUT</name></connection>
<connection>
<GID>255</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,148,130.5,179.5</points>
<connection>
<GID>260</GID>
<name>N_in1</name></connection>
<connection>
<GID>261</GID>
<name>N_in0</name></connection>
<intersection>148 6</intersection>
<intersection>170 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>130.5,170,133.5,170</points>
<connection>
<GID>257</GID>
<name>IN_1</name></connection>
<intersection>130.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>130.5,148,153,148</points>
<intersection>130.5 0</intersection>
<intersection>153 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>153,148,153,154</points>
<connection>
<GID>275</GID>
<name>IN_0</name></connection>
<intersection>148 6</intersection></vsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136.5,176,136.5,177.5</points>
<connection>
<GID>257</GID>
<name>SEL_1</name></connection>
<intersection>177.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,177.5,151.5,177.5</points>
<connection>
<GID>264</GID>
<name>N_in1</name></connection>
<connection>
<GID>268</GID>
<name>N_in0</name></connection>
<intersection>136.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137.5,176,137.5,178.5</points>
<connection>
<GID>257</GID>
<name>SEL_0</name></connection>
<intersection>178.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,178.5,151.5,178.5</points>
<connection>
<GID>265</GID>
<name>N_in1</name></connection>
<connection>
<GID>269</GID>
<name>N_in0</name></connection>
<intersection>137.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,166,141.5,168</points>
<connection>
<GID>255</GID>
<name>clock</name></connection>
<intersection>166 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>140,166,141.5,166</points>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144.5,164,144.5,165</points>
<connection>
<GID>255</GID>
<name>clear</name></connection>
<intersection>164 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>140,164,144.5,164</points>
<connection>
<GID>273</GID>
<name>IN_0</name></connection>
<intersection>144.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,158.5,138.5,161</points>
<intersection>158.5 1</intersection>
<intersection>161 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,158.5,138.5,158.5</points>
<connection>
<GID>272</GID>
<name>IN_2</name></connection>
<intersection>138.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138.5,161,139.5,161</points>
<connection>
<GID>266</GID>
<name>OUT</name></connection>
<intersection>138.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>138,156.5,139.5,156.5</points>
<connection>
<GID>272</GID>
<name>IN_1</name></connection>
<connection>
<GID>267</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,152,138.5,154.5</points>
<intersection>152 1</intersection>
<intersection>154.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138.5,152,139.5,152</points>
<connection>
<GID>270</GID>
<name>OUT</name></connection>
<intersection>138.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138,154.5,138.5,154.5</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<intersection>138.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>127,156.5,132,156.5</points>
<connection>
<GID>274</GID>
<name>N_in1</name></connection>
<connection>
<GID>272</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149.5,156.5,149.5,162</points>
<intersection>156.5 8</intersection>
<intersection>157.5 1</intersection>
<intersection>162 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145.5,157.5,149.5,157.5</points>
<connection>
<GID>267</GID>
<name>IN_1</name></connection>
<intersection>149.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>145.5,162,149.5,162</points>
<connection>
<GID>266</GID>
<name>IN_1</name></connection>
<intersection>149.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>149.5,156.5,151.5,156.5</points>
<connection>
<GID>254</GID>
<name>N_in0</name></connection>
<intersection>149.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147.5,151,147.5,160</points>
<intersection>151 3</intersection>
<intersection>154 2</intersection>
<intersection>160 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145.5,160,147.5,160</points>
<connection>
<GID>266</GID>
<name>IN_0</name></connection>
<intersection>147.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>147.5,154,149,154</points>
<connection>
<GID>275</GID>
<name>OUT_0</name></connection>
<intersection>147.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>145.5,151,147.5,151</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<intersection>147.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,149,128,174</points>
<intersection>149 2</intersection>
<intersection>174 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128,174,133.5,174</points>
<connection>
<GID>257</GID>
<name>IN_3</name></connection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>128,149,128.5,149</points>
<connection>
<GID>259</GID>
<name>N_in1</name></connection>
<intersection>128 0</intersection></hsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,172,129.5,179.5</points>
<connection>
<GID>263</GID>
<name>N_in0</name></connection>
<intersection>172 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,172,133.5,172</points>
<connection>
<GID>257</GID>
<name>IN_2</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,178.5,125,178.5</points>
<connection>
<GID>247</GID>
<name>N_in1</name></connection>
<connection>
<GID>265</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,177.5,125,177.5</points>
<connection>
<GID>246</GID>
<name>N_in1</name></connection>
<connection>
<GID>264</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,156.5,125,156.5</points>
<connection>
<GID>232</GID>
<name>N_in1</name></connection>
<connection>
<GID>274</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177,148.5,177,173.5</points>
<intersection>148.5 2</intersection>
<intersection>153 14</intersection>
<intersection>171 7</intersection>
<intersection>173.5 30</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>157,148.5,177,148.5</points>
<intersection>157 4</intersection>
<intersection>158 17</intersection>
<intersection>177 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>157,148.5,157,179.5</points>
<connection>
<GID>281</GID>
<name>N_in0</name></connection>
<intersection>148.5 2</intersection>
<intersection>168 9</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>176,171,177,171</points>
<connection>
<GID>277</GID>
<name>OUT_0</name></connection>
<intersection>177 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>157,168,162,168</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<intersection>157 4</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>174,153,177,153</points>
<connection>
<GID>293</GID>
<name>IN_1</name></connection>
<intersection>174 27</intersection>
<intersection>177 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>158,148.5,158,149</points>
<connection>
<GID>285</GID>
<name>N_in1</name></connection>
<intersection>148.5 2</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>174,153,174,155.5</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<intersection>153 14</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>170.5,173.5,177,173.5</points>
<intersection>170.5 32</intersection>
<intersection>177 0</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>170.5,173.5,170.5,175.5</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>173.5 30</intersection></vsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>168,171,170,171</points>
<connection>
<GID>279</GID>
<name>OUT</name></connection>
<connection>
<GID>277</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,148,159,179.5</points>
<connection>
<GID>283</GID>
<name>N_in1</name></connection>
<connection>
<GID>284</GID>
<name>N_in0</name></connection>
<intersection>148 6</intersection>
<intersection>170 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>159,170,162,170</points>
<connection>
<GID>279</GID>
<name>IN_1</name></connection>
<intersection>159 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>159,148,181.5,148</points>
<intersection>159 0</intersection>
<intersection>181.5 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>181.5,148,181.5,154</points>
<connection>
<GID>302</GID>
<name>IN_0</name></connection>
<intersection>148 6</intersection></vsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165,176,165,177.5</points>
<connection>
<GID>279</GID>
<name>SEL_1</name></connection>
<intersection>177.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>155.5,177.5,180,177.5</points>
<connection>
<GID>287</GID>
<name>N_in1</name></connection>
<connection>
<GID>291</GID>
<name>N_in0</name></connection>
<intersection>165 0</intersection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,176,166,178.5</points>
<connection>
<GID>279</GID>
<name>SEL_0</name></connection>
<intersection>178.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>155.5,178.5,180,178.5</points>
<connection>
<GID>288</GID>
<name>N_in1</name></connection>
<connection>
<GID>292</GID>
<name>N_in0</name></connection>
<intersection>166 0</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,166,170,168</points>
<connection>
<GID>277</GID>
<name>clock</name></connection>
<intersection>166 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168.5,166,170,166</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173,164,173,165</points>
<connection>
<GID>277</GID>
<name>clear</name></connection>
<intersection>164 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>168.5,164,173,164</points>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<intersection>173 0</intersection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,158.5,167,161</points>
<intersection>158.5 1</intersection>
<intersection>161 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166.5,158.5,167,158.5</points>
<connection>
<GID>296</GID>
<name>IN_2</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>167,161,168,161</points>
<connection>
<GID>289</GID>
<name>OUT</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>166.5,156.5,168,156.5</points>
<connection>
<GID>296</GID>
<name>IN_1</name></connection>
<connection>
<GID>290</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,152,167,154.5</points>
<intersection>152 1</intersection>
<intersection>154.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167,152,168,152</points>
<connection>
<GID>293</GID>
<name>OUT</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>166.5,154.5,167,154.5</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>155.5,156.5,160.5,156.5</points>
<connection>
<GID>300</GID>
<name>N_in1</name></connection>
<connection>
<GID>296</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178,156.5,178,162</points>
<intersection>156.5 8</intersection>
<intersection>157.5 1</intersection>
<intersection>162 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>174,157.5,178,157.5</points>
<connection>
<GID>290</GID>
<name>IN_1</name></connection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>174,162,178,162</points>
<connection>
<GID>289</GID>
<name>IN_1</name></connection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>178,156.5,180,156.5</points>
<connection>
<GID>276</GID>
<name>N_in0</name></connection>
<intersection>178 0</intersection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176,151,176,160</points>
<intersection>151 3</intersection>
<intersection>154 2</intersection>
<intersection>160 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>174,160,176,160</points>
<connection>
<GID>289</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>176,154,177.5,154</points>
<connection>
<GID>302</GID>
<name>OUT_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>174,151,176,151</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,149,156.5,174</points>
<intersection>149 2</intersection>
<intersection>174 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156.5,174,162,174</points>
<connection>
<GID>279</GID>
<name>IN_3</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156.5,149,157,149</points>
<connection>
<GID>282</GID>
<name>N_in1</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158,172,158,179.5</points>
<connection>
<GID>286</GID>
<name>N_in0</name></connection>
<intersection>172 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>158,172,162,172</points>
<connection>
<GID>279</GID>
<name>IN_2</name></connection>
<intersection>158 0</intersection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153.5,156.5,153.5,156.5</points>
<connection>
<GID>254</GID>
<name>N_in1</name></connection>
<connection>
<GID>300</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153.5,178.5,153.5,178.5</points>
<connection>
<GID>269</GID>
<name>N_in1</name></connection>
<connection>
<GID>288</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153.5,177.5,153.5,177.5</points>
<connection>
<GID>268</GID>
<name>N_in1</name></connection>
<connection>
<GID>287</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205.5,148.5,205.5,173.5</points>
<intersection>148.5 2</intersection>
<intersection>153 14</intersection>
<intersection>171 7</intersection>
<intersection>173.5 30</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>185.5,148.5,205.5,148.5</points>
<intersection>185.5 4</intersection>
<intersection>186.5 17</intersection>
<intersection>205.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>185.5,148.5,185.5,179.5</points>
<connection>
<GID>310</GID>
<name>N_in0</name></connection>
<intersection>148.5 2</intersection>
<intersection>168 9</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>204.5,171,205.5,171</points>
<connection>
<GID>306</GID>
<name>OUT_0</name></connection>
<intersection>205.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>185.5,168,190.5,168</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<intersection>185.5 4</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>202.5,153,205.5,153</points>
<connection>
<GID>223</GID>
<name>IN_1</name></connection>
<intersection>202.5 27</intersection>
<intersection>205.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>186.5,148.5,186.5,149</points>
<connection>
<GID>213</GID>
<name>N_in1</name></connection>
<intersection>148.5 2</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>202.5,153,202.5,155.5</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<intersection>153 14</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>199,173.5,205.5,173.5</points>
<intersection>199 32</intersection>
<intersection>205.5 0</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>199,173.5,199,175.5</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>173.5 30</intersection></vsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>196.5,171,198.5,171</points>
<connection>
<GID>309</GID>
<name>OUT</name></connection>
<connection>
<GID>306</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,148,187.5,179.5</points>
<connection>
<GID>312</GID>
<name>N_in1</name></connection>
<connection>
<GID>314</GID>
<name>N_in0</name></connection>
<intersection>148 6</intersection>
<intersection>170 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>187.5,170,190.5,170</points>
<connection>
<GID>309</GID>
<name>IN_1</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>187.5,148,210,148</points>
<intersection>187.5 0</intersection>
<intersection>210 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>210,148,210,154</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>148 6</intersection></vsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>193.5,176,193.5,177.5</points>
<connection>
<GID>309</GID>
<name>SEL_1</name></connection>
<intersection>177.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184,177.5,208.5,177.5</points>
<connection>
<GID>217</GID>
<name>N_in1</name></connection>
<connection>
<GID>221</GID>
<name>N_in0</name></connection>
<intersection>193.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,176,194.5,178.5</points>
<connection>
<GID>309</GID>
<name>SEL_0</name></connection>
<intersection>178.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184,178.5,208.5,178.5</points>
<connection>
<GID>218</GID>
<name>N_in1</name></connection>
<connection>
<GID>222</GID>
<name>N_in0</name></connection>
<intersection>194.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,166,198.5,168</points>
<connection>
<GID>306</GID>
<name>clock</name></connection>
<intersection>166 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>197,166,198.5,166</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201.5,164,201.5,165</points>
<connection>
<GID>306</GID>
<name>clear</name></connection>
<intersection>164 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>197,164,201.5,164</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>195.5,158.5,195.5,161</points>
<intersection>158.5 1</intersection>
<intersection>161 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>195,158.5,195.5,158.5</points>
<connection>
<GID>225</GID>
<name>IN_2</name></connection>
<intersection>195.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>195.5,161,196.5,161</points>
<connection>
<GID>219</GID>
<name>OUT</name></connection>
<intersection>195.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,156.5,196.5,156.5</points>
<connection>
<GID>225</GID>
<name>IN_1</name></connection>
<connection>
<GID>220</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>195.5,152,195.5,154.5</points>
<intersection>152 1</intersection>
<intersection>154.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>195.5,152,196.5,152</points>
<connection>
<GID>223</GID>
<name>OUT</name></connection>
<intersection>195.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>195,154.5,195.5,154.5</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>195.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>184,156.5,189,156.5</points>
<connection>
<GID>227</GID>
<name>N_in1</name></connection>
<connection>
<GID>225</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206.5,156.5,206.5,162</points>
<intersection>156.5 8</intersection>
<intersection>157.5 1</intersection>
<intersection>162 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>202.5,157.5,206.5,157.5</points>
<connection>
<GID>220</GID>
<name>IN_1</name></connection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>202.5,162,206.5,162</points>
<connection>
<GID>219</GID>
<name>IN_1</name></connection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>206.5,156.5,208.5,156.5</points>
<connection>
<GID>304</GID>
<name>N_in0</name></connection>
<intersection>206.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204.5,151,204.5,160</points>
<intersection>151 3</intersection>
<intersection>154 2</intersection>
<intersection>160 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>202.5,160,204.5,160</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>204.5,154,206,154</points>
<connection>
<GID>228</GID>
<name>OUT_0</name></connection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>202.5,151,204.5,151</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>204.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,149,185,174</points>
<intersection>149 2</intersection>
<intersection>174 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185,174,190.5,174</points>
<connection>
<GID>309</GID>
<name>IN_3</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>185,149,185.5,149</points>
<connection>
<GID>311</GID>
<name>N_in1</name></connection>
<intersection>185 0</intersection></hsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186.5,172,186.5,179.5</points>
<connection>
<GID>215</GID>
<name>N_in0</name></connection>
<intersection>172 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>186.5,172,190.5,172</points>
<connection>
<GID>309</GID>
<name>IN_2</name></connection>
<intersection>186.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182,156.5,182,156.5</points>
<connection>
<GID>227</GID>
<name>N_in0</name></connection>
<connection>
<GID>276</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182,178.5,182,178.5</points>
<connection>
<GID>218</GID>
<name>N_in0</name></connection>
<connection>
<GID>292</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182,177.5,182,177.5</points>
<connection>
<GID>217</GID>
<name>N_in0</name></connection>
<connection>
<GID>291</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210.5,156.5,210.5,156.5</points>
<connection>
<GID>230</GID>
<name>N_in0</name></connection>
<connection>
<GID>304</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211.5,157.5,211.5,179.5</points>
<connection>
<GID>230</GID>
<name>N_in3</name></connection>
<connection>
<GID>229</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211.5,149,211.5,155.5</points>
<connection>
<GID>231</GID>
<name>N_in1</name></connection>
<connection>
<GID>230</GID>
<name>N_in2</name></connection></vsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,149,80,179.5</points>
<connection>
<GID>307</GID>
<name>N_in1</name></connection>
<connection>
<GID>305</GID>
<name>N_in0</name></connection>
<intersection>172 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>80,172,81.5,172</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>80.5,156.5,94.5,156.5</points>
<connection>
<GID>303</GID>
<name>N_in0</name></connection>
<intersection>80.5 8</intersection>
<intersection>81 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>81,149,81,156.5</points>
<connection>
<GID>297</GID>
<name>N_in1</name></connection>
<intersection>156.5 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>80.5,156.5,80.5,174.5</points>
<intersection>156.5 2</intersection>
<intersection>174.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>80.5,174.5,81.5,174.5</points>
<connection>
<GID>313</GID>
<name>IN_1</name></connection>
<intersection>80.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,174,87.5,175.5</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<connection>
<GID>313</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,173,93.5,178.5</points>
<connection>
<GID>315</GID>
<name>OUT</name></connection>
<intersection>178.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93.5,178.5,94.5,178.5</points>
<connection>
<GID>299</GID>
<name>N_in0</name></connection>
<intersection>93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94.5,168,94.5,177.5</points>
<connection>
<GID>301</GID>
<name>N_in0</name></connection>
<intersection>168 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>93.5,168,94.5,168</points>
<connection>
<GID>214</GID>
<name>OUT</name></connection>
<intersection>94.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,167,81,179.5</points>
<connection>
<GID>295</GID>
<name>N_in0</name></connection>
<intersection>167 3</intersection>
<intersection>176.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81,176.5,81.5,176.5</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>81,167,87.5,167</points>
<connection>
<GID>214</GID>
<name>IN_1</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,172,88.5,172</points>
<connection>
<GID>216</GID>
<name>OUT_0</name></connection>
<connection>
<GID>315</GID>
<name>IN_1</name></connection>
<intersection>88.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>88.5,169,88.5,172</points>
<intersection>169 8</intersection>
<intersection>172 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>87.5,169,88.5,169</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>88.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,114,120,139</points>
<intersection>114 2</intersection>
<intersection>118.5 14</intersection>
<intersection>136.5 7</intersection>
<intersection>139 30</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>100,114,120,114</points>
<intersection>100 4</intersection>
<intersection>101 17</intersection>
<intersection>120 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>100,114,100,145</points>
<connection>
<GID>339</GID>
<name>N_in0</name></connection>
<intersection>114 2</intersection>
<intersection>133.5 9</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>119,136.5,120,136.5</points>
<connection>
<GID>336</GID>
<name>OUT_0</name></connection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>100,133.5,105,133.5</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<intersection>100 4</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>117,118.5,120,118.5</points>
<connection>
<GID>351</GID>
<name>IN_1</name></connection>
<intersection>117 27</intersection>
<intersection>120 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>101,114,101,114.5</points>
<connection>
<GID>343</GID>
<name>N_in1</name></connection>
<intersection>114 2</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>117,118.5,117,121</points>
<connection>
<GID>348</GID>
<name>IN_0</name></connection>
<intersection>118.5 14</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>113.5,139,120,139</points>
<intersection>113.5 32</intersection>
<intersection>120 0</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>113.5,139,113.5,141</points>
<connection>
<GID>337</GID>
<name>IN_0</name></connection>
<intersection>139 30</intersection></vsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>111,136.5,113,136.5</points>
<connection>
<GID>338</GID>
<name>OUT</name></connection>
<connection>
<GID>336</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,113.5,102,145</points>
<connection>
<GID>342</GID>
<name>N_in0</name></connection>
<connection>
<GID>341</GID>
<name>N_in1</name></connection>
<intersection>113.5 6</intersection>
<intersection>135.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>102,135.5,105,135.5</points>
<connection>
<GID>338</GID>
<name>IN_1</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>102,113.5,124.5,113.5</points>
<intersection>102 0</intersection>
<intersection>124.5 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>124.5,113.5,124.5,119.5</points>
<connection>
<GID>356</GID>
<name>IN_0</name></connection>
<intersection>113.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,141.5,108,143</points>
<connection>
<GID>338</GID>
<name>SEL_1</name></connection>
<intersection>143 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,143,123,143</points>
<connection>
<GID>349</GID>
<name>N_in0</name></connection>
<connection>
<GID>345</GID>
<name>N_in1</name></connection>
<intersection>108 0</intersection></hsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109,141.5,109,144</points>
<connection>
<GID>338</GID>
<name>SEL_0</name></connection>
<intersection>144 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,144,123,144</points>
<connection>
<GID>350</GID>
<name>N_in0</name></connection>
<connection>
<GID>346</GID>
<name>N_in1</name></connection>
<intersection>109 0</intersection></hsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,131.5,113,133.5</points>
<connection>
<GID>336</GID>
<name>clock</name></connection>
<intersection>131.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111.5,131.5,113,131.5</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<intersection>113 0</intersection></hsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,129.5,116,130.5</points>
<connection>
<GID>336</GID>
<name>clear</name></connection>
<intersection>129.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>111.5,129.5,116,129.5</points>
<connection>
<GID>354</GID>
<name>IN_0</name></connection>
<intersection>116 0</intersection></hsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,124,110,126.5</points>
<intersection>124 1</intersection>
<intersection>126.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109.5,124,110,124</points>
<connection>
<GID>353</GID>
<name>IN_2</name></connection>
<intersection>110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,126.5,111,126.5</points>
<connection>
<GID>347</GID>
<name>OUT</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109.5,122,111,122</points>
<connection>
<GID>353</GID>
<name>IN_1</name></connection>
<connection>
<GID>348</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,117.5,110,120</points>
<intersection>117.5 1</intersection>
<intersection>120 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110,117.5,111,117.5</points>
<connection>
<GID>351</GID>
<name>OUT</name></connection>
<intersection>110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109.5,120,110,120</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>98.5,122,103.5,122</points>
<connection>
<GID>355</GID>
<name>N_in1</name></connection>
<connection>
<GID>353</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,122,121,127.5</points>
<intersection>122 8</intersection>
<intersection>123 1</intersection>
<intersection>127.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117,123,121,123</points>
<connection>
<GID>348</GID>
<name>IN_1</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>117,127.5,121,127.5</points>
<connection>
<GID>347</GID>
<name>IN_1</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>121,122,123,122</points>
<connection>
<GID>335</GID>
<name>N_in0</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,116.5,119,125.5</points>
<intersection>116.5 3</intersection>
<intersection>119.5 2</intersection>
<intersection>125.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117,125.5,119,125.5</points>
<connection>
<GID>347</GID>
<name>IN_0</name></connection>
<intersection>119 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>119,119.5,120.5,119.5</points>
<connection>
<GID>356</GID>
<name>OUT_0</name></connection>
<intersection>119 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>117,116.5,119,116.5</points>
<connection>
<GID>351</GID>
<name>IN_0</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,114.5,99.5,139.5</points>
<intersection>114.5 2</intersection>
<intersection>139.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99.5,139.5,105,139.5</points>
<connection>
<GID>338</GID>
<name>IN_3</name></connection>
<intersection>99.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99.5,114.5,100,114.5</points>
<connection>
<GID>340</GID>
<name>N_in1</name></connection>
<intersection>99.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>272</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,137.5,101,145</points>
<connection>
<GID>344</GID>
<name>N_in0</name></connection>
<intersection>137.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,137.5,105,137.5</points>
<connection>
<GID>338</GID>
<name>IN_2</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>273</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,122,96.5,122</points>
<connection>
<GID>355</GID>
<name>N_in0</name></connection>
<connection>
<GID>405</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,144,96.5,144</points>
<connection>
<GID>346</GID>
<name>N_in0</name></connection>
<connection>
<GID>401</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,143,96.5,143</points>
<connection>
<GID>345</GID>
<name>N_in0</name></connection>
<connection>
<GID>403</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>276</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148.5,114,148.5,139</points>
<intersection>114 2</intersection>
<intersection>118.5 14</intersection>
<intersection>136.5 7</intersection>
<intersection>139 30</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>128.5,114,148.5,114</points>
<intersection>128.5 4</intersection>
<intersection>129.5 17</intersection>
<intersection>148.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>128.5,114,128.5,145</points>
<connection>
<GID>361</GID>
<name>N_in0</name></connection>
<intersection>114 2</intersection>
<intersection>133.5 9</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>147.5,136.5,148.5,136.5</points>
<connection>
<GID>358</GID>
<name>OUT_0</name></connection>
<intersection>148.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>128.5,133.5,133.5,133.5</points>
<connection>
<GID>360</GID>
<name>IN_0</name></connection>
<intersection>128.5 4</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>145.5,118.5,148.5,118.5</points>
<connection>
<GID>373</GID>
<name>IN_1</name></connection>
<intersection>145.5 27</intersection>
<intersection>148.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>129.5,114,129.5,114.5</points>
<connection>
<GID>365</GID>
<name>N_in1</name></connection>
<intersection>114 2</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>145.5,118.5,145.5,121</points>
<connection>
<GID>370</GID>
<name>IN_0</name></connection>
<intersection>118.5 14</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>142,139,148.5,139</points>
<intersection>142 32</intersection>
<intersection>148.5 0</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>142,139,142,141</points>
<connection>
<GID>359</GID>
<name>IN_0</name></connection>
<intersection>139 30</intersection></vsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>139.5,136.5,141.5,136.5</points>
<connection>
<GID>360</GID>
<name>OUT</name></connection>
<connection>
<GID>358</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>278</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,113.5,130.5,145</points>
<connection>
<GID>364</GID>
<name>N_in0</name></connection>
<connection>
<GID>363</GID>
<name>N_in1</name></connection>
<intersection>113.5 6</intersection>
<intersection>135.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>130.5,135.5,133.5,135.5</points>
<connection>
<GID>360</GID>
<name>IN_1</name></connection>
<intersection>130.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>130.5,113.5,153,113.5</points>
<intersection>130.5 0</intersection>
<intersection>153 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>153,113.5,153,119.5</points>
<connection>
<GID>378</GID>
<name>IN_0</name></connection>
<intersection>113.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136.5,141.5,136.5,143</points>
<connection>
<GID>360</GID>
<name>SEL_1</name></connection>
<intersection>143 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,143,151.5,143</points>
<connection>
<GID>371</GID>
<name>N_in0</name></connection>
<connection>
<GID>367</GID>
<name>N_in1</name></connection>
<intersection>136.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>280</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137.5,141.5,137.5,144</points>
<connection>
<GID>360</GID>
<name>SEL_0</name></connection>
<intersection>144 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,144,151.5,144</points>
<connection>
<GID>372</GID>
<name>N_in0</name></connection>
<connection>
<GID>368</GID>
<name>N_in1</name></connection>
<intersection>137.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>281</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,131.5,141.5,133.5</points>
<connection>
<GID>358</GID>
<name>clock</name></connection>
<intersection>131.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>140,131.5,141.5,131.5</points>
<connection>
<GID>374</GID>
<name>IN_0</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>282</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144.5,129.5,144.5,130.5</points>
<connection>
<GID>358</GID>
<name>clear</name></connection>
<intersection>129.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>140,129.5,144.5,129.5</points>
<connection>
<GID>376</GID>
<name>IN_0</name></connection>
<intersection>144.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>283</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,124,138.5,126.5</points>
<intersection>124 1</intersection>
<intersection>126.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,124,138.5,124</points>
<connection>
<GID>375</GID>
<name>IN_2</name></connection>
<intersection>138.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138.5,126.5,139.5,126.5</points>
<connection>
<GID>369</GID>
<name>OUT</name></connection>
<intersection>138.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>284</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>138,122,139.5,122</points>
<connection>
<GID>375</GID>
<name>IN_1</name></connection>
<connection>
<GID>370</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>285</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,117.5,138.5,120</points>
<intersection>117.5 1</intersection>
<intersection>120 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138.5,117.5,139.5,117.5</points>
<connection>
<GID>373</GID>
<name>OUT</name></connection>
<intersection>138.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138,120,138.5,120</points>
<connection>
<GID>375</GID>
<name>IN_0</name></connection>
<intersection>138.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>286</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>127,122,132,122</points>
<connection>
<GID>377</GID>
<name>N_in1</name></connection>
<connection>
<GID>375</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>287</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149.5,122,149.5,127.5</points>
<intersection>122 8</intersection>
<intersection>123 1</intersection>
<intersection>127.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145.5,123,149.5,123</points>
<connection>
<GID>370</GID>
<name>IN_1</name></connection>
<intersection>149.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>145.5,127.5,149.5,127.5</points>
<connection>
<GID>369</GID>
<name>IN_1</name></connection>
<intersection>149.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>149.5,122,151.5,122</points>
<connection>
<GID>357</GID>
<name>N_in0</name></connection>
<intersection>149.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>288</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147.5,116.5,147.5,125.5</points>
<intersection>116.5 3</intersection>
<intersection>119.5 2</intersection>
<intersection>125.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145.5,125.5,147.5,125.5</points>
<connection>
<GID>369</GID>
<name>IN_0</name></connection>
<intersection>147.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>147.5,119.5,149,119.5</points>
<connection>
<GID>378</GID>
<name>OUT_0</name></connection>
<intersection>147.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>145.5,116.5,147.5,116.5</points>
<connection>
<GID>373</GID>
<name>IN_0</name></connection>
<intersection>147.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>289</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,114.5,128,139.5</points>
<intersection>114.5 2</intersection>
<intersection>139.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128,139.5,133.5,139.5</points>
<connection>
<GID>360</GID>
<name>IN_3</name></connection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>128,114.5,128.5,114.5</points>
<connection>
<GID>362</GID>
<name>N_in1</name></connection>
<intersection>128 0</intersection></hsegment></shape></wire>
<wire>
<ID>290</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,137.5,129.5,145</points>
<connection>
<GID>366</GID>
<name>N_in0</name></connection>
<intersection>137.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,137.5,133.5,137.5</points>
<connection>
<GID>360</GID>
<name>IN_2</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>291</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,144,125,144</points>
<connection>
<GID>350</GID>
<name>N_in1</name></connection>
<connection>
<GID>368</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>292</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,143,125,143</points>
<connection>
<GID>349</GID>
<name>N_in1</name></connection>
<connection>
<GID>367</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>293</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,122,125,122</points>
<connection>
<GID>335</GID>
<name>N_in1</name></connection>
<connection>
<GID>377</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>294</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177,114,177,139</points>
<intersection>114 2</intersection>
<intersection>118.5 14</intersection>
<intersection>136.5 7</intersection>
<intersection>139 30</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>157,114,177,114</points>
<intersection>157 4</intersection>
<intersection>158 17</intersection>
<intersection>177 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>157,114,157,145</points>
<connection>
<GID>383</GID>
<name>N_in0</name></connection>
<intersection>114 2</intersection>
<intersection>133.5 9</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>176,136.5,177,136.5</points>
<connection>
<GID>380</GID>
<name>OUT_0</name></connection>
<intersection>177 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>157,133.5,162,133.5</points>
<connection>
<GID>382</GID>
<name>IN_0</name></connection>
<intersection>157 4</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>174,118.5,177,118.5</points>
<connection>
<GID>395</GID>
<name>IN_1</name></connection>
<intersection>174 27</intersection>
<intersection>177 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>158,114,158,114.5</points>
<connection>
<GID>387</GID>
<name>N_in1</name></connection>
<intersection>114 2</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>174,118.5,174,121</points>
<connection>
<GID>392</GID>
<name>IN_0</name></connection>
<intersection>118.5 14</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>170.5,139,177,139</points>
<intersection>170.5 32</intersection>
<intersection>177 0</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>170.5,139,170.5,141</points>
<connection>
<GID>381</GID>
<name>IN_0</name></connection>
<intersection>139 30</intersection></vsegment></shape></wire>
<wire>
<ID>295</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>168,136.5,170,136.5</points>
<connection>
<GID>382</GID>
<name>OUT</name></connection>
<connection>
<GID>380</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>296</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,113.5,159,145</points>
<connection>
<GID>386</GID>
<name>N_in0</name></connection>
<connection>
<GID>385</GID>
<name>N_in1</name></connection>
<intersection>113.5 6</intersection>
<intersection>135.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>159,135.5,162,135.5</points>
<connection>
<GID>382</GID>
<name>IN_1</name></connection>
<intersection>159 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>159,113.5,181.5,113.5</points>
<intersection>159 0</intersection>
<intersection>181.5 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>181.5,113.5,181.5,119.5</points>
<connection>
<GID>404</GID>
<name>IN_0</name></connection>
<intersection>113.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>297</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165,141.5,165,143</points>
<connection>
<GID>382</GID>
<name>SEL_1</name></connection>
<intersection>143 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>155.5,143,180,143</points>
<connection>
<GID>393</GID>
<name>N_in0</name></connection>
<connection>
<GID>389</GID>
<name>N_in1</name></connection>
<intersection>165 0</intersection></hsegment></shape></wire>
<wire>
<ID>298</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,141.5,166,144</points>
<connection>
<GID>382</GID>
<name>SEL_0</name></connection>
<intersection>144 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>155.5,144,180,144</points>
<connection>
<GID>394</GID>
<name>N_in0</name></connection>
<connection>
<GID>390</GID>
<name>N_in1</name></connection>
<intersection>166 0</intersection></hsegment></shape></wire>
<wire>
<ID>299</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,131.5,170,133.5</points>
<connection>
<GID>380</GID>
<name>clock</name></connection>
<intersection>131.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168.5,131.5,170,131.5</points>
<connection>
<GID>396</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment></shape></wire>
<wire>
<ID>300</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173,129.5,173,130.5</points>
<connection>
<GID>380</GID>
<name>clear</name></connection>
<intersection>129.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>168.5,129.5,173,129.5</points>
<connection>
<GID>400</GID>
<name>IN_0</name></connection>
<intersection>173 0</intersection></hsegment></shape></wire>
<wire>
<ID>301</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,124,167,126.5</points>
<intersection>124 1</intersection>
<intersection>126.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166.5,124,167,124</points>
<connection>
<GID>398</GID>
<name>IN_2</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>167,126.5,168,126.5</points>
<connection>
<GID>391</GID>
<name>OUT</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>302</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>166.5,122,168,122</points>
<connection>
<GID>398</GID>
<name>IN_1</name></connection>
<connection>
<GID>392</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>303</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,117.5,167,120</points>
<intersection>117.5 1</intersection>
<intersection>120 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167,117.5,168,117.5</points>
<connection>
<GID>395</GID>
<name>OUT</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>166.5,120,167,120</points>
<connection>
<GID>398</GID>
<name>IN_0</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>304</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>155.5,122,160.5,122</points>
<connection>
<GID>402</GID>
<name>N_in1</name></connection>
<connection>
<GID>398</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>305</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178,122,178,127.5</points>
<intersection>122 8</intersection>
<intersection>123 1</intersection>
<intersection>127.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>174,123,178,123</points>
<connection>
<GID>392</GID>
<name>IN_1</name></connection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>174,127.5,178,127.5</points>
<connection>
<GID>391</GID>
<name>IN_1</name></connection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>178,122,180,122</points>
<connection>
<GID>379</GID>
<name>N_in0</name></connection>
<intersection>178 0</intersection></hsegment></shape></wire>
<wire>
<ID>306</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176,116.5,176,125.5</points>
<intersection>116.5 3</intersection>
<intersection>119.5 2</intersection>
<intersection>125.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>174,125.5,176,125.5</points>
<connection>
<GID>391</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>176,119.5,177.5,119.5</points>
<connection>
<GID>404</GID>
<name>OUT_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>174,116.5,176,116.5</points>
<connection>
<GID>395</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,114.5,156.5,139.5</points>
<intersection>114.5 2</intersection>
<intersection>139.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156.5,139.5,162,139.5</points>
<connection>
<GID>382</GID>
<name>IN_3</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156.5,114.5,157,114.5</points>
<connection>
<GID>384</GID>
<name>N_in1</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>308</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158,137.5,158,145</points>
<connection>
<GID>388</GID>
<name>N_in0</name></connection>
<intersection>137.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>158,137.5,162,137.5</points>
<connection>
<GID>382</GID>
<name>IN_2</name></connection>
<intersection>158 0</intersection></hsegment></shape></wire>
<wire>
<ID>309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153.5,122,153.5,122</points>
<connection>
<GID>357</GID>
<name>N_in1</name></connection>
<connection>
<GID>402</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>310</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153.5,144,153.5,144</points>
<connection>
<GID>372</GID>
<name>N_in1</name></connection>
<connection>
<GID>390</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>311</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153.5,143,153.5,143</points>
<connection>
<GID>371</GID>
<name>N_in1</name></connection>
<connection>
<GID>389</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>312</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205.5,114,205.5,139</points>
<intersection>114 2</intersection>
<intersection>118.5 14</intersection>
<intersection>136.5 7</intersection>
<intersection>139 30</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>185.5,114,205.5,114</points>
<intersection>185.5 4</intersection>
<intersection>186.5 17</intersection>
<intersection>205.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>185.5,114,185.5,145</points>
<connection>
<GID>412</GID>
<name>N_in0</name></connection>
<intersection>114 2</intersection>
<intersection>133.5 9</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>204.5,136.5,205.5,136.5</points>
<connection>
<GID>408</GID>
<name>OUT_0</name></connection>
<intersection>205.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>185.5,133.5,190.5,133.5</points>
<connection>
<GID>411</GID>
<name>IN_0</name></connection>
<intersection>185.5 4</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>202.5,118.5,205.5,118.5</points>
<connection>
<GID>326</GID>
<name>IN_1</name></connection>
<intersection>202.5 27</intersection>
<intersection>205.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>186.5,114,186.5,114.5</points>
<connection>
<GID>316</GID>
<name>N_in1</name></connection>
<intersection>114 2</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>202.5,118.5,202.5,121</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<intersection>118.5 14</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>199,139,205.5,139</points>
<intersection>199 32</intersection>
<intersection>205.5 0</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>199,139,199,141</points>
<connection>
<GID>410</GID>
<name>IN_0</name></connection>
<intersection>139 30</intersection></vsegment></shape></wire>
<wire>
<ID>313</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>196.5,136.5,198.5,136.5</points>
<connection>
<GID>411</GID>
<name>OUT</name></connection>
<connection>
<GID>408</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>314</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,113.5,187.5,145</points>
<connection>
<GID>416</GID>
<name>N_in0</name></connection>
<connection>
<GID>414</GID>
<name>N_in1</name></connection>
<intersection>113.5 6</intersection>
<intersection>135.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>187.5,135.5,190.5,135.5</points>
<connection>
<GID>411</GID>
<name>IN_1</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>187.5,113.5,210,113.5</points>
<intersection>187.5 0</intersection>
<intersection>210 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>210,113.5,210,119.5</points>
<connection>
<GID>331</GID>
<name>IN_0</name></connection>
<intersection>113.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>315</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>193.5,141.5,193.5,143</points>
<connection>
<GID>411</GID>
<name>SEL_1</name></connection>
<intersection>143 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184,143,208.5,143</points>
<connection>
<GID>324</GID>
<name>N_in0</name></connection>
<connection>
<GID>320</GID>
<name>N_in1</name></connection>
<intersection>193.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>316</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,141.5,194.5,144</points>
<connection>
<GID>411</GID>
<name>SEL_0</name></connection>
<intersection>144 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184,144,208.5,144</points>
<connection>
<GID>325</GID>
<name>N_in0</name></connection>
<connection>
<GID>321</GID>
<name>N_in1</name></connection>
<intersection>194.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>317</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,131.5,198.5,133.5</points>
<connection>
<GID>408</GID>
<name>clock</name></connection>
<intersection>131.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>197,131.5,198.5,131.5</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<intersection>198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>318</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201.5,129.5,201.5,130.5</points>
<connection>
<GID>408</GID>
<name>clear</name></connection>
<intersection>129.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>197,129.5,201.5,129.5</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>319</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>195.5,124,195.5,126.5</points>
<intersection>124 1</intersection>
<intersection>126.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>195,124,195.5,124</points>
<connection>
<GID>328</GID>
<name>IN_2</name></connection>
<intersection>195.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>195.5,126.5,196.5,126.5</points>
<connection>
<GID>322</GID>
<name>OUT</name></connection>
<intersection>195.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>320</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,122,196.5,122</points>
<connection>
<GID>328</GID>
<name>IN_1</name></connection>
<connection>
<GID>323</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>321</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>195.5,117.5,195.5,120</points>
<intersection>117.5 1</intersection>
<intersection>120 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>195.5,117.5,196.5,117.5</points>
<connection>
<GID>326</GID>
<name>OUT</name></connection>
<intersection>195.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>195,120,195.5,120</points>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<intersection>195.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>322</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>184,122,189,122</points>
<connection>
<GID>330</GID>
<name>N_in1</name></connection>
<connection>
<GID>328</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>323</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206.5,122,206.5,127.5</points>
<intersection>122 8</intersection>
<intersection>123 1</intersection>
<intersection>127.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>202.5,123,206.5,123</points>
<connection>
<GID>323</GID>
<name>IN_1</name></connection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>202.5,127.5,206.5,127.5</points>
<connection>
<GID>322</GID>
<name>IN_1</name></connection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>206.5,122,208.5,122</points>
<connection>
<GID>406</GID>
<name>N_in0</name></connection>
<intersection>206.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>324</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204.5,116.5,204.5,125.5</points>
<intersection>116.5 3</intersection>
<intersection>119.5 2</intersection>
<intersection>125.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>202.5,125.5,204.5,125.5</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>204.5,119.5,206,119.5</points>
<connection>
<GID>331</GID>
<name>OUT_0</name></connection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>202.5,116.5,204.5,116.5</points>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<intersection>204.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>325</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,114.5,185,139.5</points>
<intersection>114.5 2</intersection>
<intersection>139.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185,139.5,190.5,139.5</points>
<connection>
<GID>411</GID>
<name>IN_3</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>185,114.5,185.5,114.5</points>
<connection>
<GID>413</GID>
<name>N_in1</name></connection>
<intersection>185 0</intersection></hsegment></shape></wire>
<wire>
<ID>326</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186.5,137.5,186.5,145</points>
<connection>
<GID>318</GID>
<name>N_in0</name></connection>
<intersection>137.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>186.5,137.5,190.5,137.5</points>
<connection>
<GID>411</GID>
<name>IN_2</name></connection>
<intersection>186.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>327</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182,122,182,122</points>
<connection>
<GID>330</GID>
<name>N_in0</name></connection>
<connection>
<GID>379</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>328</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182,144,182,144</points>
<connection>
<GID>321</GID>
<name>N_in0</name></connection>
<connection>
<GID>394</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>329</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182,143,182,143</points>
<connection>
<GID>320</GID>
<name>N_in0</name></connection>
<connection>
<GID>393</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>330</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210.5,122,210.5,122</points>
<connection>
<GID>333</GID>
<name>N_in0</name></connection>
<connection>
<GID>406</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>331</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211.5,123,211.5,145</points>
<connection>
<GID>333</GID>
<name>N_in3</name></connection>
<connection>
<GID>332</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>332</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211.5,114.5,211.5,121</points>
<connection>
<GID>334</GID>
<name>N_in1</name></connection>
<connection>
<GID>333</GID>
<name>N_in2</name></connection></vsegment></shape></wire>
<wire>
<ID>333</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,114.5,80,145</points>
<connection>
<GID>409</GID>
<name>N_in1</name></connection>
<connection>
<GID>407</GID>
<name>N_in0</name></connection>
<intersection>137.5 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>80,137.5,81.5,137.5</points>
<connection>
<GID>319</GID>
<name>IN_0</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>334</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>80.5,122,94.5,122</points>
<connection>
<GID>405</GID>
<name>N_in0</name></connection>
<intersection>80.5 8</intersection>
<intersection>81 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>81,114.5,81,122</points>
<connection>
<GID>399</GID>
<name>N_in1</name></connection>
<intersection>122 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>80.5,122,80.5,140</points>
<intersection>122 2</intersection>
<intersection>140 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>80.5,140,81.5,140</points>
<connection>
<GID>415</GID>
<name>IN_1</name></connection>
<intersection>80.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>335</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,139.5,87.5,141</points>
<connection>
<GID>417</GID>
<name>IN_0</name></connection>
<connection>
<GID>415</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>336</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,138.5,93.5,144</points>
<connection>
<GID>417</GID>
<name>OUT</name></connection>
<intersection>144 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93.5,144,94.5,144</points>
<connection>
<GID>401</GID>
<name>N_in0</name></connection>
<intersection>93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>337</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94.5,133.5,94.5,143</points>
<connection>
<GID>403</GID>
<name>N_in0</name></connection>
<intersection>133.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>93.5,133.5,94.5,133.5</points>
<connection>
<GID>317</GID>
<name>OUT</name></connection>
<intersection>94.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>338</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,132.5,81,145</points>
<connection>
<GID>397</GID>
<name>N_in0</name></connection>
<intersection>132.5 3</intersection>
<intersection>142 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81,142,81.5,142</points>
<connection>
<GID>415</GID>
<name>IN_0</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>81,132.5,87.5,132.5</points>
<connection>
<GID>317</GID>
<name>IN_1</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>339</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,137.5,87.5,137.5</points>
<connection>
<GID>417</GID>
<name>IN_1</name></connection>
<connection>
<GID>319</GID>
<name>OUT_0</name></connection>
<intersection>86.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>86.5,134.5,86.5,137.5</points>
<intersection>134.5 8</intersection>
<intersection>137.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>86.5,134.5,87.5,134.5</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<intersection>86.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>340</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,147,129.5,147</points>
<connection>
<GID>262</GID>
<name>N_in0</name></connection>
<connection>
<GID>366</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>341</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,147,130.5,147</points>
<connection>
<GID>260</GID>
<name>N_in0</name></connection>
<connection>
<GID>364</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>342</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,147,101,147</points>
<connection>
<GID>240</GID>
<name>N_in0</name></connection>
<connection>
<GID>344</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>343</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,147,102,147</points>
<connection>
<GID>238</GID>
<name>N_in0</name></connection>
<connection>
<GID>342</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>344</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,147,100,147</points>
<connection>
<GID>237</GID>
<name>N_in0</name></connection>
<connection>
<GID>339</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>345</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211.5,147,211.5,147</points>
<connection>
<GID>231</GID>
<name>N_in0</name></connection>
<connection>
<GID>332</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>346</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186.5,147,186.5,147</points>
<connection>
<GID>213</GID>
<name>N_in0</name></connection>
<connection>
<GID>318</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>347</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,147,187.5,147</points>
<connection>
<GID>312</GID>
<name>N_in0</name></connection>
<connection>
<GID>416</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>348</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185.5,147,185.5,147</points>
<connection>
<GID>311</GID>
<name>N_in0</name></connection>
<connection>
<GID>412</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>349</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,147,80,147</points>
<connection>
<GID>307</GID>
<name>N_in0</name></connection>
<connection>
<GID>407</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>350</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,147,81,147</points>
<connection>
<GID>297</GID>
<name>N_in0</name></connection>
<connection>
<GID>397</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>351</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158,147,158,147</points>
<connection>
<GID>285</GID>
<name>N_in0</name></connection>
<connection>
<GID>388</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>352</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,147,159,147</points>
<connection>
<GID>283</GID>
<name>N_in0</name></connection>
<connection>
<GID>386</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>353</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157,147,157,147</points>
<connection>
<GID>282</GID>
<name>N_in0</name></connection>
<connection>
<GID>383</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>354</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128.5,147,128.5,147</points>
<connection>
<GID>259</GID>
<name>N_in0</name></connection>
<connection>
<GID>361</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>355</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,79.5,120,104.5</points>
<intersection>79.5 2</intersection>
<intersection>84 14</intersection>
<intersection>102 7</intersection>
<intersection>104.5 30</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>100,79.5,120,79.5</points>
<intersection>100 4</intersection>
<intersection>101 17</intersection>
<intersection>120 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>100,79.5,100,110.5</points>
<connection>
<GID>441</GID>
<name>N_in0</name></connection>
<intersection>79.5 2</intersection>
<intersection>99 9</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>119,102,120,102</points>
<connection>
<GID>438</GID>
<name>OUT_0</name></connection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>100,99,105,99</points>
<connection>
<GID>440</GID>
<name>IN_0</name></connection>
<intersection>100 4</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>117,84,120,84</points>
<connection>
<GID>453</GID>
<name>IN_1</name></connection>
<intersection>117 27</intersection>
<intersection>120 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>101,79.5,101,80</points>
<connection>
<GID>445</GID>
<name>N_in1</name></connection>
<intersection>79.5 2</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>117,84,117,86.5</points>
<connection>
<GID>450</GID>
<name>IN_0</name></connection>
<intersection>84 14</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>113.5,104.5,120,104.5</points>
<intersection>113.5 32</intersection>
<intersection>120 0</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>113.5,104.5,113.5,106.5</points>
<connection>
<GID>439</GID>
<name>IN_0</name></connection>
<intersection>104.5 30</intersection></vsegment></shape></wire>
<wire>
<ID>356</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>111,102,113,102</points>
<connection>
<GID>440</GID>
<name>OUT</name></connection>
<connection>
<GID>438</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>357</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,79,102,110.5</points>
<connection>
<GID>444</GID>
<name>N_in0</name></connection>
<connection>
<GID>443</GID>
<name>N_in1</name></connection>
<intersection>79 6</intersection>
<intersection>101 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>102,101,105,101</points>
<connection>
<GID>440</GID>
<name>IN_1</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>102,79,124.5,79</points>
<intersection>102 0</intersection>
<intersection>124.5 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>124.5,79,124.5,85</points>
<connection>
<GID>458</GID>
<name>IN_0</name></connection>
<intersection>79 6</intersection></vsegment></shape></wire>
<wire>
<ID>358</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,107,108,108.5</points>
<connection>
<GID>440</GID>
<name>SEL_1</name></connection>
<intersection>108.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,108.5,123,108.5</points>
<connection>
<GID>451</GID>
<name>N_in0</name></connection>
<connection>
<GID>447</GID>
<name>N_in1</name></connection>
<intersection>108 0</intersection></hsegment></shape></wire>
<wire>
<ID>359</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109,107,109,109.5</points>
<connection>
<GID>440</GID>
<name>SEL_0</name></connection>
<intersection>109.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,109.5,123,109.5</points>
<connection>
<GID>452</GID>
<name>N_in0</name></connection>
<connection>
<GID>448</GID>
<name>N_in1</name></connection>
<intersection>109 0</intersection></hsegment></shape></wire>
<wire>
<ID>360</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,97,113,99</points>
<connection>
<GID>438</GID>
<name>clock</name></connection>
<intersection>97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111.5,97,113,97</points>
<connection>
<GID>454</GID>
<name>IN_0</name></connection>
<intersection>113 0</intersection></hsegment></shape></wire>
<wire>
<ID>361</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,95,116,96</points>
<connection>
<GID>438</GID>
<name>clear</name></connection>
<intersection>95 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>111.5,95,116,95</points>
<connection>
<GID>456</GID>
<name>IN_0</name></connection>
<intersection>116 0</intersection></hsegment></shape></wire>
<wire>
<ID>362</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,89.5,110,92</points>
<intersection>89.5 1</intersection>
<intersection>92 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109.5,89.5,110,89.5</points>
<connection>
<GID>455</GID>
<name>IN_2</name></connection>
<intersection>110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,92,111,92</points>
<connection>
<GID>449</GID>
<name>OUT</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>363</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109.5,87.5,111,87.5</points>
<connection>
<GID>455</GID>
<name>IN_1</name></connection>
<connection>
<GID>450</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>364</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,83,110,85.5</points>
<intersection>83 1</intersection>
<intersection>85.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110,83,111,83</points>
<connection>
<GID>453</GID>
<name>OUT</name></connection>
<intersection>110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109.5,85.5,110,85.5</points>
<connection>
<GID>455</GID>
<name>IN_0</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>365</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>98.5,87.5,103.5,87.5</points>
<connection>
<GID>457</GID>
<name>N_in1</name></connection>
<connection>
<GID>455</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>366</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,87.5,121,93</points>
<intersection>87.5 8</intersection>
<intersection>88.5 1</intersection>
<intersection>93 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117,88.5,121,88.5</points>
<connection>
<GID>450</GID>
<name>IN_1</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>117,93,121,93</points>
<connection>
<GID>449</GID>
<name>IN_1</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>121,87.5,123,87.5</points>
<connection>
<GID>437</GID>
<name>N_in0</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>367</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,82,119,91</points>
<intersection>82 3</intersection>
<intersection>85 2</intersection>
<intersection>91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117,91,119,91</points>
<connection>
<GID>449</GID>
<name>IN_0</name></connection>
<intersection>119 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>119,85,120.5,85</points>
<connection>
<GID>458</GID>
<name>OUT_0</name></connection>
<intersection>119 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>117,82,119,82</points>
<connection>
<GID>453</GID>
<name>IN_0</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>368</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,80,99.5,105</points>
<intersection>80 2</intersection>
<intersection>105 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99.5,105,105,105</points>
<connection>
<GID>440</GID>
<name>IN_3</name></connection>
<intersection>99.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99.5,80,100,80</points>
<connection>
<GID>442</GID>
<name>N_in1</name></connection>
<intersection>99.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>369</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,103,101,110.5</points>
<connection>
<GID>446</GID>
<name>N_in0</name></connection>
<intersection>103 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,103,105,103</points>
<connection>
<GID>440</GID>
<name>IN_2</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>370</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,87.5,96.5,87.5</points>
<connection>
<GID>457</GID>
<name>N_in0</name></connection>
<connection>
<GID>507</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>371</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,109.5,96.5,109.5</points>
<connection>
<GID>448</GID>
<name>N_in0</name></connection>
<connection>
<GID>503</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>372</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,108.5,96.5,108.5</points>
<connection>
<GID>447</GID>
<name>N_in0</name></connection>
<connection>
<GID>505</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>373</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148.5,79.5,148.5,104.5</points>
<intersection>79.5 2</intersection>
<intersection>84 14</intersection>
<intersection>102 7</intersection>
<intersection>104.5 30</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>128.5,79.5,148.5,79.5</points>
<intersection>128.5 4</intersection>
<intersection>129.5 17</intersection>
<intersection>148.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>128.5,79.5,128.5,110.5</points>
<connection>
<GID>463</GID>
<name>N_in0</name></connection>
<intersection>79.5 2</intersection>
<intersection>99 9</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>147.5,102,148.5,102</points>
<connection>
<GID>460</GID>
<name>OUT_0</name></connection>
<intersection>148.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>128.5,99,133.5,99</points>
<connection>
<GID>462</GID>
<name>IN_0</name></connection>
<intersection>128.5 4</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>145.5,84,148.5,84</points>
<connection>
<GID>475</GID>
<name>IN_1</name></connection>
<intersection>145.5 27</intersection>
<intersection>148.5 0</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>129.5,79.5,129.5,80</points>
<connection>
<GID>467</GID>
<name>N_in1</name></connection>
<intersection>79.5 2</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>145.5,84,145.5,86.5</points>
<connection>
<GID>472</GID>
<name>IN_0</name></connection>
<intersection>84 14</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>142,104.5,148.5,104.5</points>
<intersection>142 32</intersection>
<intersection>148.5 0</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>142,104.5,142,106.5</points>
<connection>
<GID>461</GID>
<name>IN_0</name></connection>
<intersection>104.5 30</intersection></vsegment></shape></wire>
<wire>
<ID>374</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>139.5,102,141.5,102</points>
<connection>
<GID>462</GID>
<name>OUT</name></connection>
<connection>
<GID>460</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>375</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,79,130.5,110.5</points>
<connection>
<GID>466</GID>
<name>N_in0</name></connection>
<connection>
<GID>465</GID>
<name>N_in1</name></connection>
<intersection>79 6</intersection>
<intersection>101 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>130.5,101,133.5,101</points>
<connection>
<GID>462</GID>
<name>IN_1</name></connection>
<intersection>130.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>130.5,79,153,79</points>
<intersection>130.5 0</intersection>
<intersection>153 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>153,79,153,85</points>
<connection>
<GID>480</GID>
<name>IN_0</name></connection>
<intersection>79 6</intersection></vsegment></shape></wire>
<wire>
<ID>376</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136.5,107,136.5,108.5</points>
<connection>
<GID>462</GID>
<name>SEL_1</name></connection>
<intersection>108.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,108.5,151.5,108.5</points>
<connection>
<GID>473</GID>
<name>N_in0</name></connection>
<connection>
<GID>469</GID>
<name>N_in1</name></connection>
<intersection>136.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>377</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137.5,107,137.5,109.5</points>
<connection>
<GID>462</GID>
<name>SEL_0</name></connection>
<intersection>109.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,109.5,151.5,109.5</points>
<connection>
<GID>474</GID>
<name>N_in0</name></connection>
<connection>
<GID>470</GID>
<name>N_in1</name></connection>
<intersection>137.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>378</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,97,141.5,99</points>
<connection>
<GID>460</GID>
<name>clock</name></connection>
<intersection>97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>140,97,141.5,97</points>
<connection>
<GID>476</GID>
<name>IN_0</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>379</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144.5,95,144.5,96</points>
<connection>
<GID>460</GID>
<name>clear</name></connection>
<intersection>95 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>140,95,144.5,95</points>
<connection>
<GID>478</GID>
<name>IN_0</name></connection>
<intersection>144.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>380</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,89.5,138.5,92</points>
<intersection>89.5 1</intersection>
<intersection>92 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,89.5,138.5,89.5</points>
<connection>
<GID>477</GID>
<name>IN_2</name></connection>
<intersection>138.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138.5,92,139.5,92</points>
<connection>
<GID>471</GID>
<name>OUT</name></connection>
<intersection>138.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>381</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>138,87.5,139.5,87.5</points>
<connection>
<GID>477</GID>
<name>IN_1</name></connection>
<connection>
<GID>472</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>382</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,83,138.5,85.5</points>
<intersection>83 1</intersection>
<intersection>85.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138.5,83,139.5,83</points>
<connection>
<GID>475</GID>
<name>OUT</name></connection>
<intersection>138.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138,85.5,138.5,85.5</points>
<connection>
<GID>477</GID>
<name>IN_0</name></connection>
<intersection>138.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>383</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>127,87.5,132,87.5</points>
<connection>
<GID>479</GID>
<name>N_in1</name></connection>
<connection>
<GID>477</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>384</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149.5,87.5,149.5,93</points>
<intersection>87.5 8</intersection>
<intersection>88.5 1</intersection>
<intersection>93 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145.5,88.5,149.5,88.5</points>
<connection>
<GID>472</GID>
<name>IN_1</name></connection>
<intersection>149.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>145.5,93,149.5,93</points>
<connection>
<GID>471</GID>
<name>IN_1</name></connection>
<intersection>149.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>149.5,87.5,151.5,87.5</points>
<connection>
<GID>459</GID>
<name>N_in0</name></connection>
<intersection>149.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>385</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147.5,82,147.5,91</points>
<intersection>82 3</intersection>
<intersection>85 2</intersection>
<intersection>91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145.5,91,147.5,91</points>
<connection>
<GID>471</GID>
<name>IN_0</name></connection>
<intersection>147.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>147.5,85,149,85</points>
<connection>
<GID>480</GID>
<name>OUT_0</name></connection>
<intersection>147.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>145.5,82,147.5,82</points>
<connection>
<GID>475</GID>
<name>IN_0</name></connection>
<intersection>147.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>386</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,80,128,105</points>
<intersection>80 2</intersection>
<intersection>105 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128,105,133.5,105</points>
<connection>
<GID>462</GID>
<name>IN_3</name></connection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>128,80,128.5,80</points>
<connection>
<GID>464</GID>
<name>N_in1</name></connection>
<intersection>128 0</intersection></hsegment></shape></wire>
<wire>
<ID>387</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,103,129.5,110.5</points>
<connection>
<GID>468</GID>
<name>N_in0</name></connection>
<intersection>103 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,103,133.5,103</points>
<connection>
<GID>462</GID>
<name>IN_2</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>388</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,109.5,125,109.5</points>
<connection>
<GID>452</GID>
<name>N_in1</name></connection>
<connection>
<GID>470</GID>
<name>N_in0</name></connection></vsegment></shape></wire></page 3>
<page 4>
<PageViewport>-98.5019,842.364,1199.5,98.3635</PageViewport></page 4>
<page 5>
<PageViewport>-98.5019,842.364,1199.5,98.3635</PageViewport></page 5>
<page 6>
<PageViewport>-98.5019,842.364,1199.5,98.3635</PageViewport></page 6>
<page 7>
<PageViewport>-98.5019,842.364,1199.5,98.3635</PageViewport></page 7>
<page 8>
<PageViewport>-98.5019,842.364,1199.5,98.3635</PageViewport></page 8>
<page 9>
<PageViewport>-98.5019,842.364,1199.5,98.3635</PageViewport></page 9></circuit>