<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-14.1687,-4.99556,102.253,-85.2501</PageViewport>
<gate>
<ID>2</ID>
<type>AA_AND2</type>
<position>72,-15</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AE_FULLADDER_4BIT</type>
<position>56,-23.5</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>34 </input>
<input>
<ID>IN_2</ID>33 </input>
<input>
<ID>IN_3</ID>32 </input>
<input>
<ID>IN_B_0</ID>39 </input>
<input>
<ID>IN_B_1</ID>38 </input>
<input>
<ID>IN_B_2</ID>37 </input>
<input>
<ID>IN_B_3</ID>36 </input>
<output>
<ID>OUT_0</ID>70 </output>
<output>
<ID>OUT_1</ID>68 </output>
<output>
<ID>OUT_2</ID>67 </output>
<output>
<ID>OUT_3</ID>66 </output>
<input>
<ID>carry_in</ID>41 </input>
<output>
<ID>carry_out</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>6</ID>
<type>DD_KEYPAD_HEX</type>
<position>16,-32</position>
<output>
<ID>OUT_0</ID>4 </output>
<output>
<ID>OUT_1</ID>3 </output>
<output>
<ID>OUT_2</ID>2 </output>
<output>
<ID>OUT_3</ID>1 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 4</lparam></gate>
<gate>
<ID>8</ID>
<type>GF_LED_DISPLAY_4BIT_OUT</type>
<position>27.5,-30</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>2 </input>
<input>
<ID>IN_3</ID>1 </input>
<output>
<ID>OUT_0</ID>8 </output>
<output>
<ID>OUT_1</ID>7 </output>
<output>
<ID>OUT_2</ID>6 </output>
<output>
<ID>OUT_3</ID>5 </output>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 4</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>10</ID>
<type>DE_TO</type>
<position>31.5,-35.5</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>11</ID>
<type>DE_TO</type>
<position>31.5,-37.5</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>12</ID>
<type>DE_TO</type>
<position>31.5,-39.5</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>13</ID>
<type>DE_TO</type>
<position>31.5,-41.5</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>14</ID>
<type>DD_KEYPAD_HEX</type>
<position>16,-49</position>
<output>
<ID>OUT_0</ID>12 </output>
<output>
<ID>OUT_1</ID>11 </output>
<output>
<ID>OUT_2</ID>10 </output>
<output>
<ID>OUT_3</ID>9 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 11</lparam></gate>
<gate>
<ID>15</ID>
<type>GF_LED_DISPLAY_4BIT_OUT</type>
<position>27.5,-47</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>11 </input>
<input>
<ID>IN_2</ID>10 </input>
<input>
<ID>IN_3</ID>9 </input>
<output>
<ID>OUT_0</ID>16 </output>
<output>
<ID>OUT_1</ID>15 </output>
<output>
<ID>OUT_2</ID>14 </output>
<output>
<ID>OUT_3</ID>13 </output>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 11</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>16</ID>
<type>DE_TO</type>
<position>31.5,-52.5</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B3</lparam></gate>
<gate>
<ID>17</ID>
<type>DE_TO</type>
<position>31.5,-54.5</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B2</lparam></gate>
<gate>
<ID>18</ID>
<type>DE_TO</type>
<position>31.5,-56.5</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B1</lparam></gate>
<gate>
<ID>19</ID>
<type>DE_TO</type>
<position>31.5,-58.5</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B0</lparam></gate>
<gate>
<ID>21</ID>
<type>DA_FROM</type>
<position>73,-8</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B0</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND2</type>
<position>68,-15</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>DA_FROM</type>
<position>69,-8</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B1</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_AND2</type>
<position>64,-15</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>DA_FROM</type>
<position>65,-8</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B2</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_AND2</type>
<position>60,-15</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>27</ID>
<type>DA_FROM</type>
<position>61,-8</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B3</lparam></gate>
<gate>
<ID>39</ID>
<type>DA_FROM</type>
<position>57.5,-8</position>
<input>
<ID>IN_0</ID>21 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_AND2</type>
<position>54,-15</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>41</ID>
<type>DA_FROM</type>
<position>55,-8</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B0</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_AND2</type>
<position>50,-15</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>43</ID>
<type>DA_FROM</type>
<position>51,-8</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B1</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_AND2</type>
<position>46,-15</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>45</ID>
<type>DA_FROM</type>
<position>47,-8</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B2</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_AND2</type>
<position>42,-15</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>DA_FROM</type>
<position>43,-8</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B3</lparam></gate>
<gate>
<ID>48</ID>
<type>DA_FROM</type>
<position>39.5,-8</position>
<input>
<ID>IN_0</ID>31 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>50</ID>
<type>FF_GND</type>
<position>57,-18.5</position>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>52</ID>
<type>HA_JUNC_2</type>
<position>72,-27</position>
<input>
<ID>N_in0</ID>69 </input>
<input>
<ID>N_in1</ID>40 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>54</ID>
<type>FF_GND</type>
<position>65,-23.5</position>
<output>
<ID>OUT_0</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>55</ID>
<type>HA_JUNC_2</type>
<position>58,-31</position>
<input>
<ID>N_in0</ID>65 </input>
<input>
<ID>N_in1</ID>42 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>57</ID>
<type>AE_FULLADDER_4BIT</type>
<position>56,-48.5</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>55 </input>
<input>
<ID>IN_2</ID>54 </input>
<input>
<ID>IN_3</ID>53 </input>
<input>
<ID>IN_B_0</ID>68 </input>
<input>
<ID>IN_B_1</ID>67 </input>
<input>
<ID>IN_B_2</ID>66 </input>
<input>
<ID>IN_B_3</ID>65 </input>
<output>
<ID>OUT_0</ID>87 </output>
<output>
<ID>OUT_1</ID>86 </output>
<output>
<ID>OUT_2</ID>85 </output>
<output>
<ID>OUT_3</ID>83 </output>
<input>
<ID>carry_in</ID>62 </input>
<output>
<ID>carry_out</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_AND2</type>
<position>54,-40</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>52 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>67</ID>
<type>DA_FROM</type>
<position>55,-33</position>
<input>
<ID>IN_0</ID>48 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B0</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_AND2</type>
<position>50,-40</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>52 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>DA_FROM</type>
<position>51,-33</position>
<input>
<ID>IN_0</ID>49 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B1</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_AND2</type>
<position>46,-40</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>52 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>71</ID>
<type>DA_FROM</type>
<position>47,-33</position>
<input>
<ID>IN_0</ID>50 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B2</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_AND2</type>
<position>42,-40</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>52 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>73</ID>
<type>DA_FROM</type>
<position>43,-33</position>
<input>
<ID>IN_0</ID>51 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B3</lparam></gate>
<gate>
<ID>74</ID>
<type>DA_FROM</type>
<position>39.5,-33</position>
<input>
<ID>IN_0</ID>52 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>76</ID>
<type>HA_JUNC_2</type>
<position>72,-75</position>
<input>
<ID>N_in0</ID>96 </input>
<input>
<ID>N_in1</ID>69 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>77</ID>
<type>FF_GND</type>
<position>65,-48.5</position>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>81</ID>
<type>HA_JUNC_2</type>
<position>71,-75</position>
<input>
<ID>N_in0</ID>95 </input>
<input>
<ID>N_in1</ID>70 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>82</ID>
<type>HA_JUNC_2</type>
<position>57.5,-56</position>
<input>
<ID>N_in0</ID>82 </input>
<input>
<ID>N_in1</ID>84 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>83</ID>
<type>AE_FULLADDER_4BIT</type>
<position>55.5,-73.5</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>78 </input>
<input>
<ID>IN_2</ID>77 </input>
<input>
<ID>IN_3</ID>76 </input>
<input>
<ID>IN_B_0</ID>86 </input>
<input>
<ID>IN_B_1</ID>85 </input>
<input>
<ID>IN_B_2</ID>83 </input>
<input>
<ID>IN_B_3</ID>82 </input>
<output>
<ID>OUT_0</ID>93 </output>
<output>
<ID>OUT_1</ID>92 </output>
<output>
<ID>OUT_2</ID>91 </output>
<output>
<ID>OUT_3</ID>90 </output>
<input>
<ID>carry_in</ID>80 </input>
<output>
<ID>carry_out</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_AND2</type>
<position>53.5,-65</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>75 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>85</ID>
<type>DA_FROM</type>
<position>54.5,-58</position>
<input>
<ID>IN_0</ID>71 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B0</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_AND2</type>
<position>49.5,-65</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>75 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>87</ID>
<type>DA_FROM</type>
<position>50.5,-58</position>
<input>
<ID>IN_0</ID>72 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B1</lparam></gate>
<gate>
<ID>88</ID>
<type>AA_AND2</type>
<position>45.5,-65</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>75 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>89</ID>
<type>DA_FROM</type>
<position>46.5,-58</position>
<input>
<ID>IN_0</ID>73 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B2</lparam></gate>
<gate>
<ID>90</ID>
<type>AA_AND2</type>
<position>41.5,-65</position>
<input>
<ID>IN_0</ID>74 </input>
<input>
<ID>IN_1</ID>75 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>91</ID>
<type>DA_FROM</type>
<position>42.5,-58</position>
<input>
<ID>IN_0</ID>74 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B3</lparam></gate>
<gate>
<ID>92</ID>
<type>DA_FROM</type>
<position>39.5,-58</position>
<input>
<ID>IN_0</ID>75 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>93</ID>
<type>FF_GND</type>
<position>64.5,-73.5</position>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>94</ID>
<type>HA_JUNC_2</type>
<position>52.5,-79</position>
<input>
<ID>N_in0</ID>89 </input>
<input>
<ID>N_in1</ID>81 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>97</ID>
<type>HA_JUNC_2</type>
<position>70,-75</position>
<input>
<ID>N_in0</ID>94 </input>
<input>
<ID>N_in1</ID>87 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>101</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>60,-82</position>
<input>
<ID>IN_0</ID>92 </input>
<input>
<ID>IN_1</ID>91 </input>
<input>
<ID>IN_2</ID>90 </input>
<input>
<ID>IN_3</ID>89 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>103</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>75.5,-82</position>
<input>
<ID>IN_0</ID>96 </input>
<input>
<ID>IN_1</ID>95 </input>
<input>
<ID>IN_2</ID>94 </input>
<input>
<ID>IN_3</ID>93 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 12</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>105</ID>
<type>AA_LABEL</type>
<position>11.5,-22.5</position>
<gparam>LABEL_TEXT 4bit Parallel Multiplier</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-29,22.5,-28</points>
<intersection>-29 1</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-29,22.5,-29</points>
<connection>
<GID>6</GID>
<name>OUT_3</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-28,24.5,-28</points>
<connection>
<GID>8</GID>
<name>IN_3</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-31,23,-29</points>
<intersection>-31 1</intersection>
<intersection>-29 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-31,23,-31</points>
<connection>
<GID>6</GID>
<name>OUT_2</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-29,24.5,-29</points>
<connection>
<GID>8</GID>
<name>IN_2</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-33,23.5,-30</points>
<intersection>-33 1</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-33,23.5,-33</points>
<connection>
<GID>6</GID>
<name>OUT_1</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23.5,-30,24.5,-30</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-35,24.5,-31</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-35,24.5,-35</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-35.5,26,-34</points>
<connection>
<GID>8</GID>
<name>OUT_3</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-35.5,29.5,-35.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-37.5,27,-34</points>
<connection>
<GID>8</GID>
<name>OUT_2</name></connection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-37.5,29.5,-37.5</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-39.5,28,-34</points>
<connection>
<GID>8</GID>
<name>OUT_1</name></connection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-39.5,29.5,-39.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-41.5,29,-34</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-41.5,29.5,-41.5</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-46,22.5,-45</points>
<intersection>-46 1</intersection>
<intersection>-45 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-46,22.5,-46</points>
<connection>
<GID>14</GID>
<name>OUT_3</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-45,24.5,-45</points>
<connection>
<GID>15</GID>
<name>IN_3</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-48,23,-46</points>
<intersection>-48 1</intersection>
<intersection>-46 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-48,23,-48</points>
<connection>
<GID>14</GID>
<name>OUT_2</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-46,24.5,-46</points>
<connection>
<GID>15</GID>
<name>IN_2</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-50,23.5,-47</points>
<intersection>-50 1</intersection>
<intersection>-47 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-50,23.5,-50</points>
<connection>
<GID>14</GID>
<name>OUT_1</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23.5,-47,24.5,-47</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-52,24.5,-48</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>-52 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-52,24.5,-52</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-52.5,26,-51</points>
<connection>
<GID>15</GID>
<name>OUT_3</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-52.5,29.5,-52.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-54.5,27,-51</points>
<connection>
<GID>15</GID>
<name>OUT_2</name></connection>
<intersection>-54.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-54.5,29.5,-54.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-56.5,28,-51</points>
<connection>
<GID>15</GID>
<name>OUT_1</name></connection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-56.5,29.5,-56.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-58.5,29,-51</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-58.5,29.5,-58.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>10</ID>
<points>73,-12,73,-10</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>21</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>9</ID>
<points>69,-12,69,-10</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<connection>
<GID>23</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>9</ID>
<points>65,-12,65,-10</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<connection>
<GID>25</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>9</ID>
<points>61,-12,61,-10</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<connection>
<GID>27</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-12,57.5,-10</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>-12 9</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-11,71,-11</points>
<intersection>57.5 0</intersection>
<intersection>63 7</intersection>
<intersection>67 6</intersection>
<intersection>71 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>71,-12,71,-11</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>-11 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>67,-12,67,-11</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>-11 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>63,-12,63,-11</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>57.5,-12,59,-12</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>10</ID>
<points>55,-12,55,-10</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<connection>
<GID>41</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>9</ID>
<points>51,-12,51,-10</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<connection>
<GID>43</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>9</ID>
<points>47,-12,47,-10</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<connection>
<GID>45</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>9</ID>
<points>43,-12,43,-10</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<connection>
<GID>47</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-12,39.5,-10</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>-12 9</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-11,53,-11</points>
<intersection>39.5 0</intersection>
<intersection>45 7</intersection>
<intersection>49 6</intersection>
<intersection>53 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>53,-12,53,-11</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>-11 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>49,-12,49,-11</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>-11 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>45,-12,45,-11</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>39.5,-12,41,-12</points>
<connection>
<GID>46</GID>
<name>IN_1</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-19.5,42,-18</points>
<connection>
<GID>46</GID>
<name>OUT</name></connection>
<intersection>-19.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>42,-19.5,51,-19.5</points>
<connection>
<GID>4</GID>
<name>IN_3</name></connection>
<intersection>42 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-19,46,-18</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>-19 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>52,-19.5,52,-19</points>
<connection>
<GID>4</GID>
<name>IN_2</name></connection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>46,-19,52,-19</points>
<intersection>46 0</intersection>
<intersection>52 1</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-19.5,53,-18.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>-18.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>50,-18.5,50,-18</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>50,-18.5,53,-18.5</points>
<intersection>50 1</intersection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-19.5,54,-18</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<connection>
<GID>40</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-19.5,58,-17.5</points>
<connection>
<GID>4</GID>
<name>IN_B_3</name></connection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>57,-17.5,58,-17.5</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>58 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-19.5,59,-18.5</points>
<connection>
<GID>4</GID>
<name>IN_B_2</name></connection>
<intersection>-18.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>60,-18.5,60,-18</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>59,-18.5,60,-18.5</points>
<intersection>59 0</intersection>
<intersection>60 1</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-19.5,60,-19</points>
<connection>
<GID>4</GID>
<name>IN_B_1</name></connection>
<intersection>-19 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>64,-19,64,-18</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>60,-19,64,-19</points>
<intersection>60 0</intersection>
<intersection>64 1</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-19.5,68,-18</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>-19.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>61,-19.5,68,-19.5</points>
<connection>
<GID>4</GID>
<name>IN_B_0</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-26,72,-18</points>
<connection>
<GID>52</GID>
<name>N_in1</name></connection>
<connection>
<GID>2</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64,-22.5,65,-22.5</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<connection>
<GID>4</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-30,47,-22.5</points>
<intersection>-30 2</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-22.5,48,-22.5</points>
<connection>
<GID>4</GID>
<name>carry_out</name></connection>
<intersection>47 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>47,-30,58,-30</points>
<connection>
<GID>55</GID>
<name>N_in1</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>10</ID>
<points>55,-37,55,-35</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<connection>
<GID>67</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>9</ID>
<points>51,-37,51,-35</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<connection>
<GID>69</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>9</ID>
<points>47,-37,47,-35</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<connection>
<GID>71</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>9</ID>
<points>43,-37,43,-35</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<connection>
<GID>73</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-37,39.5,-35</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>-37 9</intersection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-36,53,-36</points>
<intersection>39.5 0</intersection>
<intersection>45 7</intersection>
<intersection>49 6</intersection>
<intersection>53 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>53,-37,53,-36</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<intersection>-36 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>49,-37,49,-36</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<intersection>-36 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>45,-37,45,-36</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>39.5,-37,41,-37</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-44.5,42,-43</points>
<connection>
<GID>72</GID>
<name>OUT</name></connection>
<intersection>-44.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>42,-44.5,51,-44.5</points>
<connection>
<GID>57</GID>
<name>IN_3</name></connection>
<intersection>42 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-44,46,-43</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<intersection>-44 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>52,-44.5,52,-44</points>
<connection>
<GID>57</GID>
<name>IN_2</name></connection>
<intersection>-44 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>46,-44,52,-44</points>
<intersection>46 0</intersection>
<intersection>52 1</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-44.5,53,-43.5</points>
<connection>
<GID>57</GID>
<name>IN_1</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>50,-43.5,50,-43</points>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>50,-43.5,53,-43.5</points>
<intersection>50 1</intersection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-44.5,54,-43</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<connection>
<GID>66</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>64,-47.5,65,-47.5</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<connection>
<GID>57</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-44.5,58,-32</points>
<connection>
<GID>57</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>55</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-44.5,59,-29</points>
<connection>
<GID>57</GID>
<name>IN_B_2</name></connection>
<intersection>-29 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>54.5,-29,54.5,-27.5</points>
<connection>
<GID>4</GID>
<name>OUT_3</name></connection>
<intersection>-29 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>54.5,-29,59,-29</points>
<intersection>54.5 1</intersection>
<intersection>59 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-44.5,60,-28.5</points>
<connection>
<GID>57</GID>
<name>IN_B_1</name></connection>
<intersection>-28.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>55.5,-28.5,55.5,-27.5</points>
<connection>
<GID>4</GID>
<name>OUT_2</name></connection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>55.5,-28.5,60,-28.5</points>
<intersection>55.5 1</intersection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-28,56.5,-27.5</points>
<connection>
<GID>4</GID>
<name>OUT_1</name></connection>
<intersection>-28 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>61,-44.5,61,-28</points>
<connection>
<GID>57</GID>
<name>IN_B_0</name></connection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-28,61,-28</points>
<intersection>56.5 0</intersection>
<intersection>61 1</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-74,72,-28</points>
<connection>
<GID>52</GID>
<name>N_in0</name></connection>
<connection>
<GID>76</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>71,-74,71,-27.5</points>
<connection>
<GID>81</GID>
<name>N_in1</name></connection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>57.5,-27.5,71,-27.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>71 1</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>10</ID>
<points>54.5,-62,54.5,-60</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<connection>
<GID>85</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>9</ID>
<points>50.5,-62,50.5,-60</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<connection>
<GID>87</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>9</ID>
<points>46.5,-62,46.5,-60</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<connection>
<GID>89</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>9</ID>
<points>42.5,-62,42.5,-60</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<connection>
<GID>91</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-62,40.5,-60</points>
<connection>
<GID>90</GID>
<name>IN_1</name></connection>
<intersection>-61 1</intersection>
<intersection>-60 12</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-61,52.5,-61</points>
<intersection>40.5 0</intersection>
<intersection>44.5 7</intersection>
<intersection>48.5 6</intersection>
<intersection>52.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>52.5,-62,52.5,-61</points>
<connection>
<GID>84</GID>
<name>IN_1</name></connection>
<intersection>-61 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>48.5,-62,48.5,-61</points>
<connection>
<GID>86</GID>
<name>IN_1</name></connection>
<intersection>-61 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>44.5,-62,44.5,-61</points>
<connection>
<GID>88</GID>
<name>IN_1</name></connection>
<intersection>-61 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>39.5,-60,40.5,-60</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-69.5,41.5,-68</points>
<connection>
<GID>90</GID>
<name>OUT</name></connection>
<intersection>-69.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>41.5,-69.5,50.5,-69.5</points>
<connection>
<GID>83</GID>
<name>IN_3</name></connection>
<intersection>41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-69,45.5,-68</points>
<connection>
<GID>88</GID>
<name>OUT</name></connection>
<intersection>-69 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>51.5,-69.5,51.5,-69</points>
<connection>
<GID>83</GID>
<name>IN_2</name></connection>
<intersection>-69 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-69,51.5,-69</points>
<intersection>45.5 0</intersection>
<intersection>51.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-69.5,52.5,-68.5</points>
<connection>
<GID>83</GID>
<name>IN_1</name></connection>
<intersection>-68.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>49.5,-68.5,49.5,-68</points>
<connection>
<GID>86</GID>
<name>OUT</name></connection>
<intersection>-68.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-68.5,52.5,-68.5</points>
<intersection>49.5 1</intersection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-69.5,53.5,-68</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<connection>
<GID>84</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>63.5,-72.5,64.5,-72.5</points>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection>
<connection>
<GID>83</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-78,46.5,-72.5</points>
<intersection>-78 2</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-72.5,47.5,-72.5</points>
<connection>
<GID>83</GID>
<name>carry_out</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46.5,-78,52.5,-78</points>
<connection>
<GID>94</GID>
<name>N_in1</name></connection>
<intersection>46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-69.5,57.5,-57</points>
<connection>
<GID>83</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>82</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-69.5,58.5,-54.5</points>
<connection>
<GID>83</GID>
<name>IN_B_2</name></connection>
<intersection>-54.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>54.5,-54.5,54.5,-52.5</points>
<connection>
<GID>57</GID>
<name>OUT_3</name></connection>
<intersection>-54.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>54.5,-54.5,58.5,-54.5</points>
<intersection>54.5 1</intersection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-55,57.5,-55</points>
<connection>
<GID>82</GID>
<name>N_in1</name></connection>
<intersection>48 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-55,48,-47.5</points>
<connection>
<GID>57</GID>
<name>carry_out</name></connection>
<intersection>-55 1</intersection></vsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-69.5,59.5,-54</points>
<connection>
<GID>83</GID>
<name>IN_B_1</name></connection>
<intersection>-54 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>55.5,-54,55.5,-52.5</points>
<connection>
<GID>57</GID>
<name>OUT_2</name></connection>
<intersection>-54 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>55.5,-54,59.5,-54</points>
<intersection>55.5 1</intersection>
<intersection>59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-69.5,60.5,-53.5</points>
<connection>
<GID>83</GID>
<name>IN_B_0</name></connection>
<intersection>-53.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>56.5,-53.5,56.5,-52.5</points>
<connection>
<GID>57</GID>
<name>OUT_1</name></connection>
<intersection>-53.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-53.5,60.5,-53.5</points>
<intersection>56.5 1</intersection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-74,70,-52.5</points>
<connection>
<GID>97</GID>
<name>N_in1</name></connection>
<intersection>-52.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>57.5,-52.5,70,-52.5</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52.5,-80,57,-80</points>
<connection>
<GID>94</GID>
<name>N_in0</name></connection>
<connection>
<GID>101</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-81,54,-77.5</points>
<connection>
<GID>83</GID>
<name>OUT_3</name></connection>
<intersection>-81 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-81,57,-81</points>
<connection>
<GID>101</GID>
<name>IN_2</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-82,55,-77.5</points>
<connection>
<GID>83</GID>
<name>OUT_2</name></connection>
<intersection>-82 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-82,57,-82</points>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-83,56,-77.5</points>
<connection>
<GID>83</GID>
<name>OUT_1</name></connection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-83,57,-83</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-77.5,72.5,-77.5</points>
<connection>
<GID>83</GID>
<name>OUT_0</name></connection>
<intersection>72.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>72.5,-80,72.5,-77.5</points>
<connection>
<GID>103</GID>
<name>IN_3</name></connection>
<intersection>-77.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-81,70,-76</points>
<connection>
<GID>97</GID>
<name>N_in0</name></connection>
<intersection>-81 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70,-81,72.5,-81</points>
<connection>
<GID>103</GID>
<name>IN_2</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-82,71,-76</points>
<connection>
<GID>81</GID>
<name>N_in0</name></connection>
<intersection>-82 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71,-82,72.5,-82</points>
<connection>
<GID>103</GID>
<name>IN_1</name></connection>
<intersection>71 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-83,72,-76</points>
<connection>
<GID>76</GID>
<name>N_in0</name></connection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-83,72.5,-83</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-2.01941,9.79449e-007,105.619,-74.2</PageViewport></page 1>
<page 2>
<PageViewport>-2.01941,9.79449e-007,105.619,-74.2</PageViewport></page 2>
<page 3>
<PageViewport>-2.01941,9.79449e-007,105.619,-74.2</PageViewport></page 3>
<page 4>
<PageViewport>-2.01941,9.79449e-007,105.619,-74.2</PageViewport></page 4>
<page 5>
<PageViewport>-2.01941,9.79449e-007,105.619,-74.2</PageViewport></page 5>
<page 6>
<PageViewport>-2.01941,9.79449e-007,105.619,-74.2</PageViewport></page 6>
<page 7>
<PageViewport>-2.01941,9.79449e-007,105.619,-74.2</PageViewport></page 7>
<page 8>
<PageViewport>-2.01941,9.79449e-007,105.619,-74.2</PageViewport></page 8>
<page 9>
<PageViewport>-2.01941,9.79449e-007,105.619,-74.2</PageViewport></page 9></circuit>