<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>1.5,3.65194,71.9908,-52.6539</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>11.5,-11</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>11.5,-13</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>11.5,-15</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>11.5,-17</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_TOGGLE</type>
<position>8,-10</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>8,-12</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_TOGGLE</type>
<position>8,-14</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>8,-16</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AI_MUX_8x1</type>
<position>18,-13.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>8 </input>
<input>
<ID>IN_2</ID>3 </input>
<input>
<ID>IN_3</ID>7 </input>
<input>
<ID>IN_4</ID>2 </input>
<input>
<ID>IN_5</ID>6 </input>
<input>
<ID>IN_6</ID>1 </input>
<input>
<ID>IN_7</ID>5 </input>
<output>
<ID>OUT</ID>29 </output>
<input>
<ID>SEL_0</ID>168 </input>
<input>
<ID>SEL_1</ID>169 </input>
<input>
<ID>SEL_2</ID>170 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>18</ID>
<type>BB_CLOCK</type>
<position>4,-36.5</position>
<output>
<ID>CLK</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>214</ID>
<type>AA_LABEL</type>
<position>39.5,0</position>
<gparam>LABEL_TEXT Ryan Morehart</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>215</ID>
<type>AA_LABEL</type>
<position>39.5,-3.5</position>
<gparam>LABEL_TEXT Alex Laird</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AE_DFF_LOW</type>
<position>43,-13.5</position>
<input>
<ID>IN_0</ID>30 </input>
<output>
<ID>OUT_0</ID>9 </output>
<input>
<ID>clock</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>24</ID>
<type>GA_LED</type>
<position>48.5,-11.5</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AE_DFF_LOW</type>
<position>43,-23</position>
<input>
<ID>IN_0</ID>30 </input>
<output>
<ID>OUT_0</ID>10 </output>
<input>
<ID>clock</ID>22 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>26</ID>
<type>GA_LED</type>
<position>48.5,-21</position>
<input>
<ID>N_in0</ID>10 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>AE_DFF_LOW</type>
<position>43,-32.5</position>
<input>
<ID>IN_0</ID>30 </input>
<output>
<ID>OUT_0</ID>11 </output>
<input>
<ID>clock</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>28</ID>
<type>GA_LED</type>
<position>48.5,-30.5</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AE_DFF_LOW</type>
<position>43,-42</position>
<input>
<ID>IN_0</ID>30 </input>
<output>
<ID>OUT_0</ID>12 </output>
<input>
<ID>clock</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>30</ID>
<type>GA_LED</type>
<position>48.5,-40</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AE_DFF_LOW</type>
<position>61,-17.5</position>
<input>
<ID>IN_0</ID>31 </input>
<output>
<ID>OUT_0</ID>13 </output>
<input>
<ID>clock</ID>23 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>32</ID>
<type>GA_LED</type>
<position>66.5,-15.5</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AE_DFF_LOW</type>
<position>61,-27</position>
<input>
<ID>IN_0</ID>31 </input>
<output>
<ID>OUT_0</ID>14 </output>
<input>
<ID>clock</ID>21 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>66.5,-25</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AE_DFF_LOW</type>
<position>61,-36.5</position>
<input>
<ID>IN_0</ID>31 </input>
<output>
<ID>OUT_0</ID>15 </output>
<input>
<ID>clock</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>36</ID>
<type>GA_LED</type>
<position>66.5,-34.5</position>
<input>
<ID>N_in0</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AE_DFF_LOW</type>
<position>61,-46</position>
<input>
<ID>IN_0</ID>31 </input>
<output>
<ID>OUT_0</ID>16 </output>
<input>
<ID>clock</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>38</ID>
<type>GA_LED</type>
<position>66.5,-44</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>BE_DECODER_3x8</type>
<position>29.5,-36</position>
<input>
<ID>ENABLE</ID>28 </input>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>25 </input>
<input>
<ID>IN_2</ID>26 </input>
<output>
<ID>OUT_0</ID>17 </output>
<output>
<ID>OUT_1</ID>18 </output>
<output>
<ID>OUT_2</ID>19 </output>
<output>
<ID>OUT_3</ID>20 </output>
<output>
<ID>OUT_4</ID>21 </output>
<output>
<ID>OUT_5</ID>22 </output>
<output>
<ID>OUT_6</ID>23 </output>
<output>
<ID>OUT_7</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>42</ID>
<type>DA_FROM</type>
<position>23.5,-40.5</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1S0</lparam></gate>
<gate>
<ID>43</ID>
<type>DA_FROM</type>
<position>23.5,-38.5</position>
<input>
<ID>IN_0</ID>25 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1S1</lparam></gate>
<gate>
<ID>44</ID>
<type>DA_FROM</type>
<position>23.5,-36.5</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1S2</lparam></gate>
<gate>
<ID>45</ID>
<type>DA_FROM</type>
<position>14.5,-6.5</position>
<input>
<ID>IN_0</ID>168 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1S0</lparam></gate>
<gate>
<ID>46</ID>
<type>DA_FROM</type>
<position>14.5,-4.5</position>
<input>
<ID>IN_0</ID>169 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1S1</lparam></gate>
<gate>
<ID>47</ID>
<type>DA_FROM</type>
<position>14.5,-2.5</position>
<input>
<ID>IN_0</ID>170 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1S2</lparam></gate>
<gate>
<ID>49</ID>
<type>EE_VDD</type>
<position>25.5,-30.5</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>51</ID>
<type>HE_JUNC_4</type>
<position>38,-6</position>
<input>
<ID>N_in0</ID>29 </input>
<input>
<ID>N_in1</ID>31 </input>
<input>
<ID>N_in2</ID>30 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_REGISTER4</type>
<position>10.5,-30</position>
<output>
<ID>OUT_0</ID>39 </output>
<output>
<ID>OUT_1</ID>38 </output>
<output>
<ID>OUT_2</ID>37 </output>
<input>
<ID>clock</ID>35 </input>
<input>
<ID>count_enable</ID>36 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 12</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>55</ID>
<type>AA_TOGGLE</type>
<position>7,-23.5</position>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>57</ID>
<type>DE_TO</type>
<position>17.5,-28</position>
<input>
<ID>IN_0</ID>37 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1S2</lparam></gate>
<gate>
<ID>58</ID>
<type>DE_TO</type>
<position>17.5,-30</position>
<input>
<ID>IN_0</ID>38 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1S1</lparam></gate>
<gate>
<ID>59</ID>
<type>DE_TO</type>
<position>17.5,-32</position>
<input>
<ID>IN_0</ID>39 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 1S0</lparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>12,-19.5</position>
<gparam>LABEL_TEXT I0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>12,-8.5</position>
<gparam>LABEL_TEXT I6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>8.5,-7.5</position>
<gparam>LABEL_TEXT I7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>8.5,-18.5</position>
<gparam>LABEL_TEXT I1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>22.5,-12</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>49,-14</position>
<gparam>LABEL_TEXT Out7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>49,-42.5</position>
<gparam>LABEL_TEXT Out1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>67,-46.5</position>
<gparam>LABEL_TEXT Out0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>67,-18</position>
<gparam>LABEL_TEXT Out6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,-11,15,-11</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<connection>
<GID>14</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,-13,15,-13</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<connection>
<GID>14</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,-15,15,-15</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<connection>
<GID>14</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,-17,15,-17</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<connection>
<GID>14</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10,-10,15,-10</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<connection>
<GID>14</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10,-12,15,-12</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<connection>
<GID>14</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10,-14,15,-14</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<connection>
<GID>14</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10,-16,15,-16</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<connection>
<GID>14</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46,-11.5,47.5,-11.5</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<connection>
<GID>24</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46,-21,47.5,-21</points>
<connection>
<GID>26</GID>
<name>N_in0</name></connection>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46,-30.5,47.5,-30.5</points>
<connection>
<GID>28</GID>
<name>N_in0</name></connection>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46,-40,47.5,-40</points>
<connection>
<GID>30</GID>
<name>N_in0</name></connection>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64,-15.5,65.5,-15.5</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<connection>
<GID>32</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64,-25,65.5,-25</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<connection>
<GID>34</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64,-34.5,65.5,-34.5</points>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection>
<connection>
<GID>36</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64,-44,65.5,-44</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<connection>
<GID>38</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-47,33.5,-39.5</points>
<intersection>-47 1</intersection>
<intersection>-39.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-47,58,-47</points>
<connection>
<GID>37</GID>
<name>clock</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-39.5,33.5,-39.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-43,34,-38.5</points>
<intersection>-43 1</intersection>
<intersection>-38.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-43,40,-43</points>
<connection>
<GID>29</GID>
<name>clock</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-38.5,34,-38.5</points>
<connection>
<GID>40</GID>
<name>OUT_1</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32.5,-37.5,58,-37.5</points>
<connection>
<GID>35</GID>
<name>clock</name></connection>
<connection>
<GID>40</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-36.5,35,-33.5</points>
<intersection>-36.5 2</intersection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-33.5,40,-33.5</points>
<connection>
<GID>27</GID>
<name>clock</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-36.5,35,-36.5</points>
<connection>
<GID>40</GID>
<name>OUT_3</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-35.5,34.5,-28</points>
<intersection>-35.5 2</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-28,58,-28</points>
<connection>
<GID>33</GID>
<name>clock</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-35.5,34.5,-35.5</points>
<connection>
<GID>40</GID>
<name>OUT_4</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-34.5,34,-24</points>
<intersection>-34.5 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-24,40,-24</points>
<connection>
<GID>25</GID>
<name>clock</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-34.5,34,-34.5</points>
<connection>
<GID>40</GID>
<name>OUT_5</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-33.5,33.5,-18.5</points>
<intersection>-33.5 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-18.5,58,-18.5</points>
<connection>
<GID>31</GID>
<name>clock</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-33.5,33.5,-33.5</points>
<connection>
<GID>40</GID>
<name>OUT_6</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-32.5,33,-14.5</points>
<intersection>-32.5 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-14.5,40,-14.5</points>
<connection>
<GID>22</GID>
<name>clock</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-32.5,33,-32.5</points>
<connection>
<GID>40</GID>
<name>OUT_7</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-38.5,26.5,-38.5</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>26.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>26.5,-38.5,26.5,-38.5</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>-38.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-37.5,26,-36.5</points>
<intersection>-37.5 1</intersection>
<intersection>-36.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-37.5,26.5,-37.5</points>
<connection>
<GID>40</GID>
<name>IN_2</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-36.5,26,-36.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-40.5,26,-39.5</points>
<intersection>-40.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-39.5,26.5,-39.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-40.5,26,-40.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-32.5,25.5,-31.5</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-32.5,26.5,-32.5</points>
<connection>
<GID>40</GID>
<name>ENABLE</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-13.5,32.5,-6</points>
<intersection>-13.5 2</intersection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-6,37,-6</points>
<connection>
<GID>51</GID>
<name>N_in0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21,-13.5,32.5,-13.5</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-40,38,-7</points>
<connection>
<GID>51</GID>
<name>N_in2</name></connection>
<intersection>-40 1</intersection>
<intersection>-30.5 2</intersection>
<intersection>-21 3</intersection>
<intersection>-11.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-40,40,-40</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38,-30.5,40,-30.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>38,-21,40,-21</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>38,-11.5,40,-11.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-44,56,-6</points>
<intersection>-44 1</intersection>
<intersection>-34.5 3</intersection>
<intersection>-25 4</intersection>
<intersection>-15.5 5</intersection>
<intersection>-6 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-44,58,-44</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39,-6,56,-6</points>
<connection>
<GID>51</GID>
<name>N_in1</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>56,-34.5,58,-34.5</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>56,-25,58,-25</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>56,-15.5,58,-15.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-36.5,9.5,-34</points>
<connection>
<GID>53</GID>
<name>clock</name></connection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,-36.5,9.5,-36.5</points>
<connection>
<GID>18</GID>
<name>CLK</name></connection>
<intersection>9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-25,10.5,-23.5</points>
<connection>
<GID>53</GID>
<name>count_enable</name></connection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-23.5,10.5,-23.5</points>
<connection>
<GID>55</GID>
<name>OUT_0</name></connection>
<intersection>10.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-29,15,-28</points>
<intersection>-29 2</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-28,15.5,-28</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>15 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14.5,-29,15,-29</points>
<connection>
<GID>53</GID>
<name>OUT_2</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14.5,-30,15.5,-30</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>14.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>14.5,-30,14.5,-30</points>
<connection>
<GID>53</GID>
<name>OUT_1</name></connection>
<intersection>-30 1</intersection></vsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-32,15,-31</points>
<intersection>-32 1</intersection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-32,15.5,-32</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>15 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14.5,-31,15,-31</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-8,19,-6.5</points>
<connection>
<GID>14</GID>
<name>SEL_0</name></connection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16.5,-6.5,19,-6.5</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-8,18,-4.5</points>
<connection>
<GID>14</GID>
<name>SEL_1</name></connection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16.5,-4.5,18,-4.5</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-8,17,-2.5</points>
<connection>
<GID>14</GID>
<name>SEL_2</name></connection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16.5,-2.5,17,-2.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>13.1109,17.75,86.3798,-40.775</PageViewport>
<gate>
<ID>1</ID>
<type>AA_TOGGLE</type>
<position>24.5,-1.5</position>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_TOGGLE</type>
<position>24.5,-3.5</position>
<output>
<ID>OUT_0</ID>41 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_TOGGLE</type>
<position>24.5,-5.5</position>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_TOGGLE</type>
<position>24.5,-7.5</position>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_TOGGLE</type>
<position>21,-0.5</position>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_TOGGLE</type>
<position>21,-2.5</position>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>21,-4.5</position>
<output>
<ID>OUT_0</ID>46 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_TOGGLE</type>
<position>21,-6.5</position>
<output>
<ID>OUT_0</ID>47 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>212</ID>
<type>AA_LABEL</type>
<position>52.5,11</position>
<gparam>LABEL_TEXT Ryan Morehart</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AI_MUX_8x1</type>
<position>31,-4</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>47 </input>
<input>
<ID>IN_2</ID>42 </input>
<input>
<ID>IN_3</ID>46 </input>
<input>
<ID>IN_4</ID>41 </input>
<input>
<ID>IN_5</ID>45 </input>
<input>
<ID>IN_6</ID>40 </input>
<input>
<ID>IN_7</ID>44 </input>
<output>
<ID>OUT</ID>68 </output>
<input>
<ID>SEL_0</ID>84 </input>
<input>
<ID>SEL_1</ID>85 </input>
<input>
<ID>SEL_2</ID>86 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>213</ID>
<type>AA_LABEL</type>
<position>52.5,7.5</position>
<gparam>LABEL_TEXT Alex Laird</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>BB_CLOCK</type>
<position>17,-27</position>
<output>
<ID>CLK</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>21</ID>
<type>AE_DFF_LOW</type>
<position>56,-4</position>
<input>
<ID>IN_0</ID>69 </input>
<output>
<ID>OUT_0</ID>48 </output>
<input>
<ID>clock</ID>63 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>23</ID>
<type>GA_LED</type>
<position>61.5,-2</position>
<input>
<ID>N_in0</ID>48 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AE_DFF_LOW</type>
<position>56,-13.5</position>
<input>
<ID>IN_0</ID>69 </input>
<output>
<ID>OUT_0</ID>49 </output>
<input>
<ID>clock</ID>61 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>41</ID>
<type>GA_LED</type>
<position>61.5,-11.5</position>
<input>
<ID>N_in0</ID>49 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AE_DFF_LOW</type>
<position>56,-23</position>
<input>
<ID>IN_0</ID>69 </input>
<output>
<ID>OUT_0</ID>50 </output>
<input>
<ID>clock</ID>59 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>50</ID>
<type>GA_LED</type>
<position>61.5,-21</position>
<input>
<ID>N_in0</ID>50 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AE_DFF_LOW</type>
<position>56,-32.5</position>
<input>
<ID>IN_0</ID>69 </input>
<output>
<ID>OUT_0</ID>51 </output>
<input>
<ID>clock</ID>57 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>54</ID>
<type>GA_LED</type>
<position>61.5,-30.5</position>
<input>
<ID>N_in0</ID>51 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AE_DFF_LOW</type>
<position>74,-8</position>
<input>
<ID>IN_0</ID>70 </input>
<output>
<ID>OUT_0</ID>52 </output>
<input>
<ID>clock</ID>62 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>60</ID>
<type>GA_LED</type>
<position>79.5,-6</position>
<input>
<ID>N_in0</ID>52 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AE_DFF_LOW</type>
<position>74,-17.5</position>
<input>
<ID>IN_0</ID>70 </input>
<output>
<ID>OUT_0</ID>53 </output>
<input>
<ID>clock</ID>60 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>71</ID>
<type>GA_LED</type>
<position>79.5,-15.5</position>
<input>
<ID>N_in0</ID>53 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>AE_DFF_LOW</type>
<position>74,-27</position>
<input>
<ID>IN_0</ID>70 </input>
<output>
<ID>OUT_0</ID>54 </output>
<input>
<ID>clock</ID>58 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>73</ID>
<type>GA_LED</type>
<position>79.5,-25</position>
<input>
<ID>N_in0</ID>54 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>AE_DFF_LOW</type>
<position>74,-36.5</position>
<input>
<ID>IN_0</ID>70 </input>
<output>
<ID>OUT_0</ID>55 </output>
<input>
<ID>clock</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>75</ID>
<type>GA_LED</type>
<position>79.5,-34.5</position>
<input>
<ID>N_in0</ID>55 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>BE_DECODER_3x8</type>
<position>42.5,-26.5</position>
<input>
<ID>ENABLE</ID>67 </input>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_1</ID>64 </input>
<input>
<ID>IN_2</ID>65 </input>
<output>
<ID>OUT_0</ID>56 </output>
<output>
<ID>OUT_1</ID>57 </output>
<output>
<ID>OUT_2</ID>58 </output>
<output>
<ID>OUT_3</ID>59 </output>
<output>
<ID>OUT_4</ID>60 </output>
<output>
<ID>OUT_5</ID>61 </output>
<output>
<ID>OUT_6</ID>62 </output>
<output>
<ID>OUT_7</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>77</ID>
<type>DA_FROM</type>
<position>36.5,-31</position>
<input>
<ID>IN_0</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 2S0</lparam></gate>
<gate>
<ID>78</ID>
<type>DA_FROM</type>
<position>36.5,-29</position>
<input>
<ID>IN_0</ID>64 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 2S1</lparam></gate>
<gate>
<ID>79</ID>
<type>DA_FROM</type>
<position>36.5,-27</position>
<input>
<ID>IN_0</ID>65 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 2S2</lparam></gate>
<gate>
<ID>83</ID>
<type>EE_VDD</type>
<position>38.5,-21</position>
<output>
<ID>OUT_0</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>84</ID>
<type>HE_JUNC_4</type>
<position>51,3.5</position>
<input>
<ID>N_in0</ID>68 </input>
<input>
<ID>N_in1</ID>70 </input>
<input>
<ID>N_in2</ID>69 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>AA_REGISTER4</type>
<position>23.5,-20.5</position>
<output>
<ID>OUT_0</ID>78 </output>
<output>
<ID>OUT_1</ID>77 </output>
<output>
<ID>OUT_2</ID>76 </output>
<input>
<ID>clock</ID>74 </input>
<input>
<ID>count_enable</ID>75 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 12</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_TOGGLE</type>
<position>20,-14</position>
<output>
<ID>OUT_0</ID>75 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>87</ID>
<type>DE_TO</type>
<position>30.5,-18.5</position>
<input>
<ID>IN_0</ID>76 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 2S2</lparam></gate>
<gate>
<ID>88</ID>
<type>DE_TO</type>
<position>30.5,-20.5</position>
<input>
<ID>IN_0</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 2S1</lparam></gate>
<gate>
<ID>89</ID>
<type>DE_TO</type>
<position>30.5,-22.5</position>
<input>
<ID>IN_0</ID>78 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 2S0</lparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>25,-10</position>
<gparam>LABEL_TEXT I0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>25,1</position>
<gparam>LABEL_TEXT I6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>AA_LABEL</type>
<position>21.5,2</position>
<gparam>LABEL_TEXT I7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>93</ID>
<type>AA_LABEL</type>
<position>21.5,-9</position>
<gparam>LABEL_TEXT I1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>94</ID>
<type>AA_LABEL</type>
<position>35.5,-2.5</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>95</ID>
<type>AA_LABEL</type>
<position>62,-4.5</position>
<gparam>LABEL_TEXT Out7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>AA_LABEL</type>
<position>62,-33</position>
<gparam>LABEL_TEXT Out1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>97</ID>
<type>AA_LABEL</type>
<position>80,-37</position>
<gparam>LABEL_TEXT Out0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>98</ID>
<type>AA_LABEL</type>
<position>80,-8.5</position>
<gparam>LABEL_TEXT Out6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>100</ID>
<type>DD_KEYPAD_HEX</type>
<position>22,11.5</position>
<output>
<ID>OUT_0</ID>84 </output>
<output>
<ID>OUT_1</ID>85 </output>
<output>
<ID>OUT_2</ID>86 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-1.5,28,-1.5</points>
<connection>
<GID>19</GID>
<name>IN_6</name></connection>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-3.5,28,-3.5</points>
<connection>
<GID>19</GID>
<name>IN_4</name></connection>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-5.5,28,-5.5</points>
<connection>
<GID>19</GID>
<name>IN_2</name></connection>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-7.5,28,-7.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23,-0.5,28,-0.5</points>
<connection>
<GID>19</GID>
<name>IN_7</name></connection>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23,-2.5,28,-2.5</points>
<connection>
<GID>19</GID>
<name>IN_5</name></connection>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23,-4.5,28,-4.5</points>
<connection>
<GID>19</GID>
<name>IN_3</name></connection>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23,-6.5,28,-6.5</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59,-2,60.5,-2</points>
<connection>
<GID>23</GID>
<name>N_in0</name></connection>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59,-11.5,60.5,-11.5</points>
<connection>
<GID>41</GID>
<name>N_in0</name></connection>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59,-21,60.5,-21</points>
<connection>
<GID>50</GID>
<name>N_in0</name></connection>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59,-30.5,60.5,-30.5</points>
<connection>
<GID>54</GID>
<name>N_in0</name></connection>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>77,-6,78.5,-6</points>
<connection>
<GID>60</GID>
<name>N_in0</name></connection>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>77,-15.5,78.5,-15.5</points>
<connection>
<GID>71</GID>
<name>N_in0</name></connection>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>77,-25,78.5,-25</points>
<connection>
<GID>73</GID>
<name>N_in0</name></connection>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>77,-34.5,78.5,-34.5</points>
<connection>
<GID>75</GID>
<name>N_in0</name></connection>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-37.5,46.5,-30</points>
<intersection>-37.5 1</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-37.5,71,-37.5</points>
<connection>
<GID>74</GID>
<name>clock</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-30,46.5,-30</points>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection>
<intersection>46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-33.5,47,-29</points>
<intersection>-33.5 1</intersection>
<intersection>-29 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-33.5,53,-33.5</points>
<connection>
<GID>52</GID>
<name>clock</name></connection>
<intersection>47 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-29,47,-29</points>
<connection>
<GID>76</GID>
<name>OUT_1</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-28,71,-28</points>
<connection>
<GID>76</GID>
<name>OUT_2</name></connection>
<connection>
<GID>72</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-27,48,-24</points>
<intersection>-27 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-24,53,-24</points>
<connection>
<GID>48</GID>
<name>clock</name></connection>
<intersection>48 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-27,48,-27</points>
<connection>
<GID>76</GID>
<name>OUT_3</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-26,47.5,-18.5</points>
<intersection>-26 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-18.5,71,-18.5</points>
<connection>
<GID>70</GID>
<name>clock</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-26,47.5,-26</points>
<connection>
<GID>76</GID>
<name>OUT_4</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-25,47,-14.5</points>
<intersection>-25 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-14.5,53,-14.5</points>
<connection>
<GID>39</GID>
<name>clock</name></connection>
<intersection>47 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-25,47,-25</points>
<connection>
<GID>76</GID>
<name>OUT_5</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-24,46.5,-9</points>
<intersection>-24 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-9,71,-9</points>
<connection>
<GID>56</GID>
<name>clock</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-24,46.5,-24</points>
<connection>
<GID>76</GID>
<name>OUT_6</name></connection>
<intersection>46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-23,46,-5</points>
<intersection>-23 2</intersection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-5,53,-5</points>
<connection>
<GID>21</GID>
<name>clock</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-23,46,-23</points>
<connection>
<GID>76</GID>
<name>OUT_7</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38.5,-29,39.5,-29</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>39.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>39.5,-29,39.5,-29</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>-29 1</intersection></vsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-28,39,-27</points>
<intersection>-28 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-28,39.5,-28</points>
<connection>
<GID>76</GID>
<name>IN_2</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38.5,-27,39,-27</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-31,39,-30</points>
<intersection>-31 2</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-30,39.5,-30</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38.5,-31,39,-31</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-23,38.5,-22</points>
<connection>
<GID>83</GID>
<name>OUT_0</name></connection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-23,39.5,-23</points>
<connection>
<GID>76</GID>
<name>ENABLE</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-4,45.5,3.5</points>
<intersection>-4 2</intersection>
<intersection>3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45.5,3.5,50,3.5</points>
<connection>
<GID>84</GID>
<name>N_in0</name></connection>
<intersection>45.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-4,45.5,-4</points>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<intersection>45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-30.5,51,2.5</points>
<connection>
<GID>84</GID>
<name>N_in2</name></connection>
<intersection>-30.5 1</intersection>
<intersection>-21 2</intersection>
<intersection>-11.5 3</intersection>
<intersection>-2 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-30.5,53,-30.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51,-21,53,-21</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>51,-11.5,53,-11.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>51,-2,53,-2</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-34.5,69,3.5</points>
<intersection>-34.5 1</intersection>
<intersection>-25 3</intersection>
<intersection>-15.5 4</intersection>
<intersection>-6 5</intersection>
<intersection>3.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69,-34.5,71,-34.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>69 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,3.5,69,3.5</points>
<connection>
<GID>84</GID>
<name>N_in1</name></connection>
<intersection>69 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>69,-25,71,-25</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>69 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>69,-15.5,71,-15.5</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>69 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>69,-6,71,-6</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-27,22.5,-24.5</points>
<connection>
<GID>85</GID>
<name>clock</name></connection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-27,22.5,-27</points>
<connection>
<GID>20</GID>
<name>CLK</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-15.5,23.5,-14</points>
<connection>
<GID>85</GID>
<name>count_enable</name></connection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-14,23.5,-14</points>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-19.5,28,-18.5</points>
<intersection>-19.5 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-18.5,28.5,-18.5</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-19.5,28,-19.5</points>
<connection>
<GID>85</GID>
<name>OUT_2</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-20.5,28.5,-20.5</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>27.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>27.5,-20.5,27.5,-20.5</points>
<connection>
<GID>85</GID>
<name>OUT_1</name></connection>
<intersection>-20.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-22.5,28,-21.5</points>
<intersection>-22.5 1</intersection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-22.5,28.5,-22.5</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-21.5,28,-21.5</points>
<connection>
<GID>85</GID>
<name>OUT_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,1.5,32,8.5</points>
<connection>
<GID>19</GID>
<name>SEL_0</name></connection>
<intersection>8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,8.5,32,8.5</points>
<connection>
<GID>100</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,1.5,31,10.5</points>
<connection>
<GID>19</GID>
<name>SEL_1</name></connection>
<intersection>10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,10.5,31,10.5</points>
<connection>
<GID>100</GID>
<name>OUT_1</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,1.5,30,12.5</points>
<connection>
<GID>19</GID>
<name>SEL_2</name></connection>
<intersection>12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,12.5,30,12.5</points>
<connection>
<GID>100</GID>
<name>OUT_2</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>15.5,4.65194,85.9908,-51.6539</PageViewport>
<gate>
<ID>193</ID>
<type>AA_LABEL</type>
<position>63,-13</position>
<gparam>LABEL_TEXT Out7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>194</ID>
<type>AA_LABEL</type>
<position>63,-41.5</position>
<gparam>LABEL_TEXT Out1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>195</ID>
<type>AA_LABEL</type>
<position>81,-45.5</position>
<gparam>LABEL_TEXT Out0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>196</ID>
<type>AA_LABEL</type>
<position>81,-17</position>
<gparam>LABEL_TEXT Out6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>206</ID>
<type>AE_SMALL_INVERTER</type>
<position>37,-35.5</position>
<input>
<ID>IN_0</ID>180 </input>
<output>
<ID>OUT_0</ID>181 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>207</ID>
<type>AE_SMALL_INVERTER</type>
<position>37,-37.5</position>
<input>
<ID>IN_0</ID>183 </input>
<output>
<ID>OUT_0</ID>184 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>208</ID>
<type>AE_SMALL_INVERTER</type>
<position>37,-39.5</position>
<input>
<ID>IN_0</ID>182 </input>
<output>
<ID>OUT_0</ID>185 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>210</ID>
<type>AA_LABEL</type>
<position>52.5,1</position>
<gparam>LABEL_TEXT Ryan Morehart</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>211</ID>
<type>AA_LABEL</type>
<position>52.5,-2.5</position>
<gparam>LABEL_TEXT Alex Laird</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>148</ID>
<type>AA_TOGGLE</type>
<position>25.5,-10</position>
<output>
<ID>OUT_0</ID>126 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>149</ID>
<type>AA_TOGGLE</type>
<position>25.5,-12</position>
<output>
<ID>OUT_0</ID>127 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>150</ID>
<type>AA_TOGGLE</type>
<position>25.5,-14</position>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_TOGGLE</type>
<position>25.5,-16</position>
<output>
<ID>OUT_0</ID>129 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>152</ID>
<type>AA_TOGGLE</type>
<position>22,-9</position>
<output>
<ID>OUT_0</ID>130 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_TOGGLE</type>
<position>22,-11</position>
<output>
<ID>OUT_0</ID>131 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>154</ID>
<type>AA_TOGGLE</type>
<position>22,-13</position>
<output>
<ID>OUT_0</ID>132 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>155</ID>
<type>AA_TOGGLE</type>
<position>22,-15</position>
<output>
<ID>OUT_0</ID>133 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>156</ID>
<type>AI_MUX_8x1</type>
<position>32,-12.5</position>
<input>
<ID>IN_0</ID>129 </input>
<input>
<ID>IN_1</ID>133 </input>
<input>
<ID>IN_2</ID>128 </input>
<input>
<ID>IN_3</ID>132 </input>
<input>
<ID>IN_4</ID>127 </input>
<input>
<ID>IN_5</ID>131 </input>
<input>
<ID>IN_6</ID>126 </input>
<input>
<ID>IN_7</ID>130 </input>
<output>
<ID>OUT</ID>154 </output>
<input>
<ID>SEL_0</ID>171 </input>
<input>
<ID>SEL_1</ID>172 </input>
<input>
<ID>SEL_2</ID>173 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>157</ID>
<type>BB_CLOCK</type>
<position>18,-35.5</position>
<output>
<ID>CLK</ID>160 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>158</ID>
<type>AE_DFF_LOW</type>
<position>57,-12.5</position>
<input>
<ID>IN_0</ID>155 </input>
<output>
<ID>OUT_0</ID>134 </output>
<input>
<ID>clock</ID>149 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>159</ID>
<type>GA_LED</type>
<position>62.5,-10.5</position>
<input>
<ID>N_in0</ID>134 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>160</ID>
<type>AE_DFF_LOW</type>
<position>57,-22</position>
<input>
<ID>IN_0</ID>155 </input>
<output>
<ID>OUT_0</ID>135 </output>
<input>
<ID>clock</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>161</ID>
<type>GA_LED</type>
<position>62.5,-20</position>
<input>
<ID>N_in0</ID>135 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>162</ID>
<type>AE_DFF_LOW</type>
<position>57,-31.5</position>
<input>
<ID>IN_0</ID>155 </input>
<output>
<ID>OUT_0</ID>136 </output>
<input>
<ID>clock</ID>145 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>163</ID>
<type>GA_LED</type>
<position>62.5,-29.5</position>
<input>
<ID>N_in0</ID>136 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>164</ID>
<type>AE_DFF_LOW</type>
<position>57,-41</position>
<input>
<ID>IN_0</ID>155 </input>
<output>
<ID>OUT_0</ID>137 </output>
<input>
<ID>clock</ID>143 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>165</ID>
<type>GA_LED</type>
<position>62.5,-39</position>
<input>
<ID>N_in0</ID>137 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>166</ID>
<type>AE_DFF_LOW</type>
<position>75,-16.5</position>
<input>
<ID>IN_0</ID>156 </input>
<output>
<ID>OUT_0</ID>138 </output>
<input>
<ID>clock</ID>148 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>167</ID>
<type>GA_LED</type>
<position>80.5,-14.5</position>
<input>
<ID>N_in0</ID>138 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>168</ID>
<type>AE_DFF_LOW</type>
<position>75,-26</position>
<input>
<ID>IN_0</ID>156 </input>
<output>
<ID>OUT_0</ID>139 </output>
<input>
<ID>clock</ID>146 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>169</ID>
<type>GA_LED</type>
<position>80.5,-24</position>
<input>
<ID>N_in0</ID>139 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>AE_DFF_LOW</type>
<position>75,-35.5</position>
<input>
<ID>IN_0</ID>156 </input>
<output>
<ID>OUT_0</ID>140 </output>
<input>
<ID>clock</ID>144 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>171</ID>
<type>GA_LED</type>
<position>80.5,-33.5</position>
<input>
<ID>N_in0</ID>140 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>172</ID>
<type>AE_DFF_LOW</type>
<position>75,-45</position>
<input>
<ID>IN_0</ID>156 </input>
<output>
<ID>OUT_0</ID>141 </output>
<input>
<ID>clock</ID>142 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>173</ID>
<type>GA_LED</type>
<position>80.5,-43</position>
<input>
<ID>N_in0</ID>141 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>174</ID>
<type>BE_DECODER_3x8</type>
<position>43.5,-35</position>
<input>
<ID>ENABLE</ID>153 </input>
<input>
<ID>IN_0</ID>185 </input>
<input>
<ID>IN_1</ID>184 </input>
<input>
<ID>IN_2</ID>181 </input>
<output>
<ID>OUT_0</ID>142 </output>
<output>
<ID>OUT_1</ID>143 </output>
<output>
<ID>OUT_2</ID>144 </output>
<output>
<ID>OUT_3</ID>145 </output>
<output>
<ID>OUT_4</ID>146 </output>
<output>
<ID>OUT_5</ID>147 </output>
<output>
<ID>OUT_6</ID>148 </output>
<output>
<ID>OUT_7</ID>149 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>175</ID>
<type>DA_FROM</type>
<position>32,-39.5</position>
<input>
<ID>IN_0</ID>182 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 3S0</lparam></gate>
<gate>
<ID>176</ID>
<type>DA_FROM</type>
<position>32,-37.5</position>
<input>
<ID>IN_0</ID>183 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 3S1</lparam></gate>
<gate>
<ID>177</ID>
<type>DA_FROM</type>
<position>32,-35.5</position>
<input>
<ID>IN_0</ID>180 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 3S2</lparam></gate>
<gate>
<ID>178</ID>
<type>DA_FROM</type>
<position>28.5,-5.5</position>
<input>
<ID>IN_0</ID>171 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 3S0</lparam></gate>
<gate>
<ID>179</ID>
<type>DA_FROM</type>
<position>28.5,-3.5</position>
<input>
<ID>IN_0</ID>172 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 3S1</lparam></gate>
<gate>
<ID>180</ID>
<type>DA_FROM</type>
<position>28.5,-1.5</position>
<input>
<ID>IN_0</ID>173 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 3S2</lparam></gate>
<gate>
<ID>181</ID>
<type>EE_VDD</type>
<position>39.5,-29.5</position>
<output>
<ID>OUT_0</ID>153 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>182</ID>
<type>HE_JUNC_4</type>
<position>52,-5</position>
<input>
<ID>N_in0</ID>154 </input>
<input>
<ID>N_in1</ID>156 </input>
<input>
<ID>N_in2</ID>155 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>183</ID>
<type>AA_REGISTER4</type>
<position>24.5,-29</position>
<output>
<ID>OUT_0</ID>164 </output>
<output>
<ID>OUT_1</ID>163 </output>
<output>
<ID>OUT_2</ID>162 </output>
<input>
<ID>clock</ID>160 </input>
<input>
<ID>count_enable</ID>161 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>184</ID>
<type>AA_TOGGLE</type>
<position>21,-22.5</position>
<output>
<ID>OUT_0</ID>161 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>185</ID>
<type>DE_TO</type>
<position>31.5,-27</position>
<input>
<ID>IN_0</ID>162 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 3S2</lparam></gate>
<gate>
<ID>186</ID>
<type>DE_TO</type>
<position>31.5,-29</position>
<input>
<ID>IN_0</ID>163 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 3S1</lparam></gate>
<gate>
<ID>187</ID>
<type>DE_TO</type>
<position>31.5,-31</position>
<input>
<ID>IN_0</ID>164 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID 3S0</lparam></gate>
<gate>
<ID>188</ID>
<type>AA_LABEL</type>
<position>26,-18.5</position>
<gparam>LABEL_TEXT I0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>189</ID>
<type>AA_LABEL</type>
<position>26,-7.5</position>
<gparam>LABEL_TEXT I6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>190</ID>
<type>AA_LABEL</type>
<position>22.5,-6.5</position>
<gparam>LABEL_TEXT I7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>191</ID>
<type>AA_LABEL</type>
<position>22.5,-17.5</position>
<gparam>LABEL_TEXT I1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>192</ID>
<type>AA_LABEL</type>
<position>36.5,-11</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>126</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-10,29,-10</points>
<connection>
<GID>156</GID>
<name>IN_6</name></connection>
<connection>
<GID>148</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-12,29,-12</points>
<connection>
<GID>156</GID>
<name>IN_4</name></connection>
<connection>
<GID>149</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-14,29,-14</points>
<connection>
<GID>156</GID>
<name>IN_2</name></connection>
<connection>
<GID>150</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-16,29,-16</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-9,29,-9</points>
<connection>
<GID>156</GID>
<name>IN_7</name></connection>
<connection>
<GID>152</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-11,29,-11</points>
<connection>
<GID>156</GID>
<name>IN_5</name></connection>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-13,29,-13</points>
<connection>
<GID>156</GID>
<name>IN_3</name></connection>
<connection>
<GID>154</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-15,29,-15</points>
<connection>
<GID>156</GID>
<name>IN_1</name></connection>
<connection>
<GID>155</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-10.5,61.5,-10.5</points>
<connection>
<GID>159</GID>
<name>N_in0</name></connection>
<connection>
<GID>158</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-20,61.5,-20</points>
<connection>
<GID>161</GID>
<name>N_in0</name></connection>
<connection>
<GID>160</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-29.5,61.5,-29.5</points>
<connection>
<GID>163</GID>
<name>N_in0</name></connection>
<connection>
<GID>162</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-39,61.5,-39</points>
<connection>
<GID>165</GID>
<name>N_in0</name></connection>
<connection>
<GID>164</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-14.5,79.5,-14.5</points>
<connection>
<GID>167</GID>
<name>N_in0</name></connection>
<connection>
<GID>166</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-24,79.5,-24</points>
<connection>
<GID>169</GID>
<name>N_in0</name></connection>
<connection>
<GID>168</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-33.5,79.5,-33.5</points>
<connection>
<GID>171</GID>
<name>N_in0</name></connection>
<connection>
<GID>170</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-43,79.5,-43</points>
<connection>
<GID>173</GID>
<name>N_in0</name></connection>
<connection>
<GID>172</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-46,47.5,-38.5</points>
<intersection>-46 1</intersection>
<intersection>-38.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-46,72,-46</points>
<connection>
<GID>172</GID>
<name>clock</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46.5,-38.5,47.5,-38.5</points>
<connection>
<GID>174</GID>
<name>OUT_0</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-42,48,-37.5</points>
<intersection>-42 1</intersection>
<intersection>-37.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-42,54,-42</points>
<connection>
<GID>164</GID>
<name>clock</name></connection>
<intersection>48 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46.5,-37.5,48,-37.5</points>
<connection>
<GID>174</GID>
<name>OUT_1</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-36.5,72,-36.5</points>
<connection>
<GID>174</GID>
<name>OUT_2</name></connection>
<connection>
<GID>170</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-35.5,49,-32.5</points>
<intersection>-35.5 2</intersection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-32.5,54,-32.5</points>
<connection>
<GID>162</GID>
<name>clock</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46.5,-35.5,49,-35.5</points>
<connection>
<GID>174</GID>
<name>OUT_3</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,-34.5,48.5,-27</points>
<intersection>-34.5 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48.5,-27,72,-27</points>
<connection>
<GID>168</GID>
<name>clock</name></connection>
<intersection>48.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46.5,-34.5,48.5,-34.5</points>
<connection>
<GID>174</GID>
<name>OUT_4</name></connection>
<intersection>48.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-33.5,48,-23</points>
<intersection>-33.5 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-23,54,-23</points>
<connection>
<GID>160</GID>
<name>clock</name></connection>
<intersection>48 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46.5,-33.5,48,-33.5</points>
<connection>
<GID>174</GID>
<name>OUT_5</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-32.5,47.5,-17.5</points>
<intersection>-32.5 2</intersection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-17.5,72,-17.5</points>
<connection>
<GID>166</GID>
<name>clock</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46.5,-32.5,47.5,-32.5</points>
<connection>
<GID>174</GID>
<name>OUT_6</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-31.5,47,-13.5</points>
<intersection>-31.5 2</intersection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-13.5,54,-13.5</points>
<connection>
<GID>158</GID>
<name>clock</name></connection>
<intersection>47 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46.5,-31.5,47,-31.5</points>
<connection>
<GID>174</GID>
<name>OUT_7</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-31.5,39.5,-30.5</points>
<connection>
<GID>181</GID>
<name>OUT_0</name></connection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-31.5,40.5,-31.5</points>
<connection>
<GID>174</GID>
<name>ENABLE</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-12.5,46.5,-5</points>
<intersection>-12.5 2</intersection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-5,51,-5</points>
<connection>
<GID>182</GID>
<name>N_in0</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-12.5,46.5,-12.5</points>
<connection>
<GID>156</GID>
<name>OUT</name></connection>
<intersection>46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-39,52,-6</points>
<connection>
<GID>182</GID>
<name>N_in2</name></connection>
<intersection>-39 1</intersection>
<intersection>-29.5 2</intersection>
<intersection>-20 3</intersection>
<intersection>-10.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-39,54,-39</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,-29.5,54,-29.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>52,-20,54,-20</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>52,-10.5,54,-10.5</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-43,70,-5</points>
<intersection>-43 1</intersection>
<intersection>-33.5 3</intersection>
<intersection>-24 4</intersection>
<intersection>-14.5 5</intersection>
<intersection>-5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70,-43,72,-43</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>70 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53,-5,70,-5</points>
<connection>
<GID>182</GID>
<name>N_in1</name></connection>
<intersection>70 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>70,-33.5,72,-33.5</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>70 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>70,-24,72,-24</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>70 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>70,-14.5,72,-14.5</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-35.5,23.5,-33</points>
<connection>
<GID>183</GID>
<name>clock</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-35.5,23.5,-35.5</points>
<connection>
<GID>157</GID>
<name>CLK</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-24,24.5,-22.5</points>
<connection>
<GID>183</GID>
<name>count_enable</name></connection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-22.5,24.5,-22.5</points>
<connection>
<GID>184</GID>
<name>OUT_0</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-28,29,-27</points>
<intersection>-28 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-27,29.5,-27</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-28,29,-28</points>
<connection>
<GID>183</GID>
<name>OUT_2</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-29,29.5,-29</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>28.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>28.5,-29,28.5,-29</points>
<connection>
<GID>183</GID>
<name>OUT_1</name></connection>
<intersection>-29 1</intersection></vsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-31,29,-30</points>
<intersection>-31 1</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-31,29.5,-31</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-30,29,-30</points>
<connection>
<GID>183</GID>
<name>OUT_0</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-7,33,-5.5</points>
<connection>
<GID>156</GID>
<name>SEL_0</name></connection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-5.5,33,-5.5</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-7,32,-3.5</points>
<connection>
<GID>156</GID>
<name>SEL_1</name></connection>
<intersection>-3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-3.5,32,-3.5</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-7,31,-1.5</points>
<connection>
<GID>156</GID>
<name>SEL_2</name></connection>
<intersection>-1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-1.5,31,-1.5</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-35.5,35,-35.5</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<connection>
<GID>206</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-36.5,39.5,-35.5</points>
<intersection>-36.5 1</intersection>
<intersection>-35.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-36.5,40.5,-36.5</points>
<connection>
<GID>174</GID>
<name>IN_2</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39,-35.5,39.5,-35.5</points>
<connection>
<GID>206</GID>
<name>OUT_0</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-39.5,35,-39.5</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<connection>
<GID>175</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-37.5,35,-37.5</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<connection>
<GID>176</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39,-37.5,40.5,-37.5</points>
<connection>
<GID>207</GID>
<name>OUT_0</name></connection>
<connection>
<GID>174</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-39.5,39.5,-38.5</points>
<intersection>-39.5 2</intersection>
<intersection>-38.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-38.5,40.5,-38.5</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39,-39.5,39.5,-39.5</points>
<connection>
<GID>208</GID>
<name>OUT_0</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>0,17.3876,287.788,-212.488</PageViewport></page 3>
<page 4>
<PageViewport>0,17.3876,287.788,-212.488</PageViewport></page 4>
<page 5>
<PageViewport>0,17.3876,287.788,-212.488</PageViewport></page 5>
<page 6>
<PageViewport>0,17.3876,287.788,-212.488</PageViewport></page 6>
<page 7>
<PageViewport>0,17.3876,287.788,-212.488</PageViewport></page 7>
<page 8>
<PageViewport>0,17.3876,287.788,-212.488</PageViewport></page 8>
<page 9>
<PageViewport>0,17.3876,287.788,-212.488</PageViewport></page 9></circuit>