<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>0,0,129.8,-74.4</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>6.5,-5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>6.5,-8</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>6.5,-11</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>DE_TO</type>
<position>12.5,-5</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>10</ID>
<type>DE_TO</type>
<position>12.5,-8</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>12</ID>
<type>DE_TO</type>
<position>12.5,-11</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>14</ID>
<type>DA_FROM</type>
<position>24.5,-6</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>16</ID>
<type>DA_FROM</type>
<position>24.5,-8</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>20</ID>
<type>AI_XOR2</type>
<position>31.5,-7</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AI_XOR2</type>
<position>40.5,-8</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>DA_FROM</type>
<position>32.5,-11</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>26</ID>
<type>DE_TO</type>
<position>45.5,-8</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum</lparam></gate>
<gate>
<ID>28</ID>
<type>DA_FROM</type>
<position>61.5,-7</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Carry</lparam></gate>
<gate>
<ID>30</ID>
<type>DA_FROM</type>
<position>61.5,-9</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Sum</lparam></gate>
<gate>
<ID>32</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>68.5,-7</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>9 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>34</ID>
<type>DA_FROM</type>
<position>24.5,-16</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>36</ID>
<type>DA_FROM</type>
<position>24.5,-18</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_AND2</type>
<position>31,-17</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_AND2</type>
<position>31,-22</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_AND2</type>
<position>31,-27</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>46</ID>
<type>AE_OR2</type>
<position>39.5,-21</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>AE_OR2</type>
<position>47.5,-26</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>DA_FROM</type>
<position>24.5,-21</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>52</ID>
<type>DA_FROM</type>
<position>24.5,-23</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>54</ID>
<type>DA_FROM</type>
<position>24.5,-26</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>56</ID>
<type>DA_FROM</type>
<position>24.5,-28</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>58</ID>
<type>DE_TO</type>
<position>52.5,-26</position>
<input>
<ID>IN_0</ID>22 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Carry</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8.5,-5,10.5,-5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>8.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>8.5,-5,8.5,-5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8.5,-8,10.5,-8</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>8.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>8.5,-8,8.5,-8</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-8 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8.5,-11,10.5,-11</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>8.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>8.5,-11,8.5,-11</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>-11 1</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-6,28.5,-6</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<connection>
<GID>20</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-8,28.5,-8</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<connection>
<GID>20</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34.5,-7,37.5,-7</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<connection>
<GID>22</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-11,36,-9</points>
<intersection>-11 1</intersection>
<intersection>-9 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-11,36,-11</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36,-9,37.5,-9</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-8,43.5,-8</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-8,43.5,-8</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>63.5,-7,65.5,-7</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<connection>
<GID>32</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-9,64.5,-8</points>
<intersection>-9 2</intersection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64.5,-8,65.5,-8</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-9,64.5,-9</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-16,28,-16</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<connection>
<GID>38</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-18,28,-18</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<connection>
<GID>38</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-21,28,-21</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<connection>
<GID>50</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-23,28,-23</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<connection>
<GID>52</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-26,28,-26</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<connection>
<GID>54</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-28,28,-28</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<connection>
<GID>56</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-20,35,-17</points>
<intersection>-20 4</intersection>
<intersection>-17 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>35,-20,36.5,-20</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>34,-17,35,-17</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-22,36.5,-22</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<connection>
<GID>46</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-25,43.5,-21</points>
<intersection>-25 4</intersection>
<intersection>-21 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>43.5,-25,44.5,-25</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>42.5,-21,43.5,-21</points>
<connection>
<GID>46</GID>
<name>OUT</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-27,44.5,-27</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<connection>
<GID>48</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-26,50.5,-26</points>
<connection>
<GID>48</GID>
<name>OUT</name></connection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-26,50.5,-26</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,129.8,-74.4</PageViewport></page 1>
<page 2>
<PageViewport>0,0,129.8,-74.4</PageViewport></page 2>
<page 3>
<PageViewport>0,0,129.8,-74.4</PageViewport></page 3>
<page 4>
<PageViewport>0,0,129.8,-74.4</PageViewport></page 4>
<page 5>
<PageViewport>0,0,129.8,-74.4</PageViewport></page 5>
<page 6>
<PageViewport>0,0,129.8,-74.4</PageViewport></page 6>
<page 7>
<PageViewport>0,0,129.8,-74.4</PageViewport></page 7>
<page 8>
<PageViewport>0,0,129.8,-74.4</PageViewport></page 8>
<page 9>
<PageViewport>0,0,129.8,-74.4</PageViewport></page 9></circuit>